
`timescale 1ns/100ps

module dff (q, d,clk);

input clk, d;
output q;
reg q;
always @(posedge clk) 
q = d;

endmodule

// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND58

module c499 (PNN1,PNN5,PNN9,PNN13,PNN17,PNN21,PNN25,PNN29,PNN33,PNN37,
             PNN41,PNN45,PNN49,PNN53,PNN57,PNN61,PNN65,PNN69,PNN73,PNN77,
             PNN81,PNN85,PNN89,PNN93,PNN97,PNN101,PNN105,PNN109,PNN113,PNN117,
             PNN121,PNN125,PNN129,PNN130,PNN131,PNN132,PNN133,PNN134,PNN135,PNN136,
             PNN137,PNN724,PNN725,PNN726,PNN727,PNN728,PNN729,PNN730,PNN731,PNN732,
             PNN733,PNN734,PNN735,PNN736,PNN737,PNN738,PNN739,PNN740,PNN741,PNN742,
             PNN743,PNN744,PNN745,PNN746,PNN747,PNN748,PNN749,PNN750,PNN751,PNN752,
             PNN753,PNN754,PNN755);

input PNN1,PNN5,PNN9,PNN13,PNN17,PNN21,PNN25,PNN29,PNN33,PNN37,
      PNN41,PNN45,PNN49,PNN53,PNN57,PNN61,PNN65,PNN69,PNN73,PNN77,
      PNN81,PNN85,PNN89,PNN93,PNN97,PNN101,PNN105,PNN109,PNN113,PNN117,
      PNN121,PNN125,PNN129,PNN130,PNN131,PNN132,PNN133,PNN134,PNN135,PNN136,
      PNN137;

output PNN724,PNN725,PNN726,PNN727,PNN728,PNN729,PNN730,PNN731,PNN732,PNN733,
       PNN734,PNN735,PNN736,PNN737,PNN738,PNN739,PNN740,PNN741,PNN742,PNN743,
       PNN744,PNN745,PNN746,PNN747,PNN748,PNN749,PNN750,PNN751,PNN752,PNN753,
       PNN754,PNN755;

wire PNN250,PNN251,PNN252,PNN253,PNN254,PNN255,PNN256,PNN257,PNN258,PNN259,
     PNN260,PNN261,PNN262,PNN263,PNN264,PNN265,PNN266,PNN267,PNN268,PNN269,
     PNN270,PNN271,PNN272,PNN273,PNN274,PNN275,PNN276,PNN277,PNN278,PNN279,
     PNN280,PNN281,PNN282,PNN283,PNN284,PNN285,PNN286,PNN287,PNN288,PNN289,
     PNN290,PNN293,PNN296,PNN299,PNN302,PNN305,PNN308,PNN311,PNN314,PNN315,
     PNN316,PNN317,PNN318,PNN319,PNN320,PNN321,PNN338,PNN339,PNN340,PNN341,
     PNN342,PNN343,PNN344,PNN345,PNN346,PNN347,PNN348,PNN349,PNN350,PNN351,
     PNN352,PNN353,PNN354,PNN367,PNN380,PNN393,PNN406,PNN419,PNN432,PNN445,
     PNN554,PNN555,PNN556,PNN557,PNN558,PNN559,PNN560,PNN561,PNN562,PNN563,
     PNN564,PNN565,PNN566,PNN567,PNN568,PNN569,PNN570,PNN571,PNN572,PNN573,
     PNN574,PNN575,PNN576,PNN577,PNN578,PNN579,PNN580,PNN581,PNN582,PNN583,
     PNN584,PNN585,PNN586,PNN587,PNN588,PNN589,PNN590,PNN591,PNN592,PNN593,
     PNN594,PNN595,PNN596,PNN597,PNN598,PNN599,PNN600,PNN601,PNN602,PNN607,
     PNN620,PNN625,PNN630,PNN635,PNN640,PNN645,PNN650,PNN655,PNN692,PNN693,
     PNN694,PNN695,PNN696,PNN697,PNN698,PNN699,PNN700,PNN701,PNN702,PNN703,
     PNN704,PNN705,PNN706,PNN707,PNN708,PNN709,PNN710,PNN711,PNN712,PNN713,
     PNN714,PNN715,PNN716,PNN717,PNN718,PNN719,PNN720,PNN721,PNN722,PNN723;

xor XOR2_1 (PNN250, PNN1, PNN5);
xor XOR2_2 (PNN251, PNN9, PNN13);
xor XOR2_3 (PNN252, PNN17, PNN21);
xor XOR2_4 (PNN253, PNN25, PNN29);
xor XOR2_5 (PNN254, PNN33, PNN37);
xor XOR2_6 (PNN255, PNN41, PNN45);
xor XOR2_7 (PNN256, PNN49, PNN53);
xor XOR2_8 (PNN257, PNN57, PNN61);
xor XOR2_9 (PNN258, PNN65, PNN69);
xor XOR2_10 (PNN259, PNN73, PNN77);
xor XOR2_11 (PNN260, PNN81, PNN85);
xor XOR2_12 (PNN261, PNN89, PNN93);
xor XOR2_13 (PNN262, PNN97, PNN101);
xor XOR2_14 (PNN263, PNN105, PNN109);
xor XOR2_15 (PNN264, PNN113, PNN117);
xor XOR2_16 (PNN265, PNN121, PNN125);
and AND2_17 (PNN266, PNN129, PNN137);
and AND2_18 (PNN267, PNN130, PNN137);
and AND2_19 (PNN268, PNN131, PNN137);
and AND2_20 (PNN269, PNN132, PNN137);
and AND2_21 (PNN270, PNN133, PNN137);
and AND2_22 (PNN271, PNN134, PNN137);
and AND2_23 (PNN272, PNN135, PNN137);
and AND2_24 (PNN273, PNN136, PNN137);
xor XOR2_25 (PNN274, PNN1, PNN17);
xor XOR2_26 (PNN275, PNN33, PNN49);
xor XOR2_27 (PNN276, PNN5, PNN21);
xor XOR2_28 (PNN277, PNN37, PNN53);
xor XOR2_29 (PNN278, PNN9, PNN25);
xor XOR2_30 (PNN279, PNN41, PNN57);
xor XOR2_31 (PNN280, PNN13, PNN29);
xor XOR2_32 (PNN281, PNN45, PNN61);
xor XOR2_33 (PNN282, PNN65, PNN81);
xor XOR2_34 (PNN283, PNN97, PNN113);
xor XOR2_35 (PNN284, PNN69, PNN85);
xor XOR2_36 (PNN285, PNN101, PNN117);
xor XOR2_37 (PNN286, PNN73, PNN89);
xor XOR2_38 (PNN287, PNN105, PNN121);
xor XOR2_39 (PNN288, PNN77, PNN93);
xor XOR2_40 (PNN289, PNN109, PNN125);
xor XOR2_41 (PNN290, PNN250, PNN251);
xor XOR2_42 (PNN293, PNN252, PNN253);
xor XOR2_43 (PNN296, PNN254, PNN255);
xor XOR2_44 (PNN299, PNN256, PNN257);
xor XOR2_45 (PNN302, PNN258, PNN259);
xor XOR2_46 (PNN305, PNN260, PNN261);
xor XOR2_47 (PNN308, PNN262, PNN263);
xor XOR2_48 (PNN311, PNN264, PNN265);
xor XOR2_49 (PNN314, PNN274, PNN275);
xor XOR2_50 (PNN315, PNN276, PNN277);
xor XOR2_51 (PNN316, PNN278, PNN279);
xor XOR2_52 (PNN317, PNN280, PNN281);
xor XOR2_53 (PNN318, PNN282, PNN283);
xor XOR2_54 (PNN319, PNN284, PNN285);
xor XOR2_55 (PNN320, PNN286, PNN287);
xor XOR2_56 (PNN321, PNN288, PNN289);
xor XOR2_57 (PNN338, PNN290, PNN293);
xor XOR2_58 (PNN339, PNN296, PNN299);
xor XOR2_59 (PNN340, PNN290, PNN296);
xor XOR2_60 (PNN341, PNN293, PNN299);
xor XOR2_61 (PNN342, PNN302, PNN305);
xor XOR2_62 (PNN343, PNN308, PNN311);
xor XOR2_63 (PNN344, PNN302, PNN308);
xor XOR2_64 (PNN345, PNN305, PNN311);
xor XOR2_65 (PNN346, PNN266, PNN342);
xor XOR2_66 (PNN347, PNN267, PNN343);
xor XOR2_67 (PNN348, PNN268, PNN344);
xor XOR2_68 (PNN349, PNN269, PNN345);
xor XOR2_69 (PNN350, PNN270, PNN338);
xor XOR2_70 (PNN351, PNN271, PNN339);
xor XOR2_71 (PNN352, PNN272, PNN340);
xor XOR2_72 (PNN353, PNN273, PNN341);
xor XOR2_73 (PNN354, PNN314, PNN346);
xor XOR2_74 (PNN367, PNN315, PNN347);
xor XOR2_75 (PNN380, PNN316, PNN348);
xor XOR2_76 (PNN393, PNN317, PNN349);
xor XOR2_77 (PNN406, PNN318, PNN350);
xor XOR2_78 (PNN419, PNN319, PNN351);
xor XOR2_79 (PNN432, PNN320, PNN352);
xor XOR2_80 (PNN445, PNN321, PNN353);
not NOT1_81 (PNN554, PNN354);
not NOT1_82 (PNN555, PNN367);
not NOT1_83 (PNN556, PNN380);
not NOT1_84 (PNN557, PNN354);
not NOT1_85 (PNN558, PNN367);
not NOT1_86 (PNN559, PNN393);
not NOT1_87 (PNN560, PNN354);
not NOT1_88 (PNN561, PNN380);
not NOT1_89 (PNN562, PNN393);
not NOT1_90 (PNN563, PNN367);
not NOT1_91 (PNN564, PNN380);
not NOT1_92 (PNN565, PNN393);
not NOT1_93 (PNN566, PNN419);
not NOT1_94 (PNN567, PNN445);
not NOT1_95 (PNN568, PNN419);
not NOT1_96 (PNN569, PNN432);
not NOT1_97 (PNN570, PNN406);
not NOT1_98 (PNN571, PNN445);
not NOT1_99 (PNN572, PNN406);
not NOT1_100 (PNN573, PNN432);
not NOT1_101 (PNN574, PNN406);
not NOT1_102 (PNN575, PNN419);
not NOT1_103 (PNN576, PNN432);
not NOT1_104 (PNN577, PNN406);
not NOT1_105 (PNN578, PNN419);
not NOT1_106 (PNN579, PNN445);
not NOT1_107 (PNN580, PNN406);
not NOT1_108 (PNN581, PNN432);
not NOT1_109 (PNN582, PNN445);
not NOT1_110 (PNN583, PNN419);
not NOT1_111 (PNN584, PNN432);
not NOT1_112 (PNN585, PNN445);
not NOT1_113 (PNN586, PNN367);
not NOT1_114 (PNN587, PNN393);
not NOT1_115 (PNN588, PNN367);
not NOT1_116 (PNN589, PNN380);
not NOT1_117 (PNN590, PNN354);
not NOT1_118 (PNN591, PNN393);
not NOT1_119 (PNN592, PNN354);
not NOT1_120 (PNN593, PNN380);
and AND4_121 (PNN594, PNN554, PNN555, PNN556, PNN393);
and AND4_122 (PNN595, PNN557, PNN558, PNN380, PNN559);
and AND4_123 (PNN596, PNN560, PNN367, PNN561, PNN562);
and AND4_124 (PNN597, PNN354, PNN563, PNN564, PNN565);
and AND4_125 (PNN598, PNN574, PNN575, PNN576, PNN445);
and AND4_126 (PNN599, PNN577, PNN578, PNN432, PNN579);
and AND4_127 (PNN600, PNN580, PNN419, PNN581, PNN582);
and AND4_128 (PNN601, PNN406, PNN583, PNN584, PNN585);
or OR4_129 (PNN602, PNN594, PNN595, PNN596, PNN597);
or OR4_130 (PNN607, PNN598, PNN599, PNN600, PNN601);
and APNND5_131 (PNN620, PNN406, PNN566, PNN432, PNN567, PNN602);
and APNND5_132 (PNN625, PNN406, PNN568, PNN569, PNN445, PNN602);
and APNND5_133 (PNN630, PNN570, PNN419, PNN432, PNN571, PNN602);
and APNND5_134 (PNN635, PNN572, PNN419, PNN573, PNN445, PNN602);
and APNND5_135 (PNN640, PNN354, PNN586, PNN380, PNN587, PNN607);
and APNND5_136 (PNN645, PNN354, PNN588, PNN589, PNN393, PNN607);
and APNND5_137 (PNN650, PNN590, PNN367, PNN380, PNN591, PNN607);
and APNND5_138 (PNN655, PNN592, PNN367, PNN593, PNN393, PNN607);
and AND2_139 (PNN692, PNN354, PNN620);
and AND2_140 (PNN693, PNN367, PNN620);
and AND2_141 (PNN694, PNN380, PNN620);
and AND2_142 (PNN695, PNN393, PNN620);
and AND2_143 (PNN696, PNN354, PNN625);
and AND2_144 (PNN697, PNN367, PNN625);
and AND2_145 (PNN698, PNN380, PNN625);
and AND2_146 (PNN699, PNN393, PNN625);
and AND2_147 (PNN700, PNN354, PNN630);
and AND2_148 (PNN701, PNN367, PNN630);
and AND2_149 (PNN702, PNN380, PNN630);
and AND2_150 (PNN703, PNN393, PNN630);
and AND2_151 (PNN704, PNN354, PNN635);
and AND2_152 (PNN705, PNN367, PNN635);
and AND2_153 (PNN706, PNN380, PNN635);
and AND2_154 (PNN707, PNN393, PNN635);
and AND2_155 (PNN708, PNN406, PNN640);
and AND2_156 (PNN709, PNN419, PNN640);
and AND2_157 (PNN710, PNN432, PNN640);
and AND2_158 (PNN711, PNN445, PNN640);
and AND2_159 (PNN712, PNN406, PNN645);
and AND2_160 (PNN713, PNN419, PNN645);
and AND2_161 (PNN714, PNN432, PNN645);
and AND2_162 (PNN715, PNN445, PNN645);
and AND2_163 (PNN716, PNN406, PNN650);
and AND2_164 (PNN717, PNN419, PNN650);
and AND2_165 (PNN718, PNN432, PNN650);
and AND2_166 (PNN719, PNN445, PNN650);
and AND2_167 (PNN720, PNN406, PNN655);
and AND2_168 (PNN721, PNN419, PNN655);
and AND2_169 (PNN722, PNN432, PNN655);
and AND2_170 (PNN723, PNN445, PNN655);
xor XOR2_171 (PNN724, PNN1, PNN692);
xor XOR2_172 (PNN725, PNN5, PNN693);
xor XOR2_173 (PNN726, PNN9, PNN694);
xor XOR2_174 (PNN727, PNN13, PNN695);
xor XOR2_175 (PNN728, PNN17, PNN696);
xor XOR2_176 (PNN729, PNN21, PNN697);
xor XOR2_177 (PNN730, PNN25, PNN698);
xor XOR2_178 (PNN731, PNN29, PNN699);
xor XOR2_179 (PNN732, PNN33, PNN700);
xor XOR2_180 (PNN733, PNN37, PNN701);
xor XOR2_181 (PNN734, PNN41, PNN702);
xor XOR2_182 (PNN735, PNN45, PNN703);
xor XOR2_183 (PNN736, PNN49, PNN704);
xor XOR2_184 (PNN737, PNN53, PNN705);
xor XOR2_185 (PNN738, PNN57, PNN706);
xor XOR2_186 (PNN739, PNN61, PNN707);
xor XOR2_187 (PNN740, PNN65, PNN708);
xor XOR2_188 (PNN741, PNN69, PNN709);
xor XOR2_189 (PNN742, PNN73, PNN710);
xor XOR2_190 (PNN743, PNN77, PNN711);
xor XOR2_191 (PNN744, PNN81, PNN712);
xor XOR2_192 (PNN745, PNN85, PNN713);
xor XOR2_193 (PNN746, PNN89, PNN714);
xor XOR2_194 (PNN747, PNN93, PNN715);
xor XOR2_195 (PNN748, PNN97, PNN716);
xor XOR2_196 (PNN749, PNN101, PNN717);
xor XOR2_197 (PNN750, PNN105, PNN718);
xor XOR2_198 (PNN751, PNN109, PNN719);
xor XOR2_199 (PNN752, PNN113, PNN720);
xor XOR2_200 (PNN753, PNN117, PNN721);
xor XOR2_201 (PNN754, PNN121, PNN722);
xor XOR2_202 (PNN755, PNN125, PNN723);

endmodule



module c499_clk_ipFF (clk,PNN1,PNN5,PNN9,PNN13,PNN17,PNN21,PNN25,PNN29,PNN33,PNN37,
             PNN41,PNN45,PNN49,PNN53,PNN57,PNN61,PNN65,PNN69,PNN73,PNN77,
             PNN81,PNN85,PNN89,PNN93,PNN97,PNN101,PNN105,PNN109,PNN113,PNN117,
             PNN121,PNN125,PNN129,PNN130,PNN131,PNN132,PNN133,PNN134,PNN135,PNN136,
             PNN137,
	     Q_PNN724,Q_PNN725,Q_PNN726,Q_PNN727,Q_PNN728,Q_PNN729,Q_PNN730,Q_PNN731,Q_PNN732,
             Q_PNN733,Q_PNN734,Q_PNN735,Q_PNN736,Q_PNN737,Q_PNN738,Q_PNN739,Q_PNN740,Q_PNN741,Q_PNN742,
             Q_PNN743,Q_PNN744,Q_PNN745,Q_PNN746,Q_PNN747,Q_PNN748,Q_PNN749,Q_PNN750,Q_PNN751,Q_PNN752,
             Q_PNN753,Q_PNN754,Q_PNN755);

input clk,PNN1,PNN5,PNN9,PNN13,PNN17,PNN21,PNN25,PNN29,PNN33,PNN37,
      PNN41,PNN45,PNN49,PNN53,PNN57,PNN61,PNN65,PNN69,PNN73,PNN77,
      PNN81,PNN85,PNN89,PNN93,PNN97,PNN101,PNN105,PNN109,PNN113,PNN117,
      PNN121,PNN125,PNN129,PNN130,PNN131,PNN132,PNN133,PNN134,PNN135,PNN136,
      PNN137;

output  Q_PNN724,Q_PNN725,Q_PNN726,Q_PNN727,Q_PNN728,Q_PNN729,Q_PNN730,Q_PNN731,Q_PNN732,
             Q_PNN733,Q_PNN734,Q_PNN735,Q_PNN736,Q_PNN737,Q_PNN738,Q_PNN739,Q_PNN740,Q_PNN741,Q_PNN742,
             Q_PNN743,Q_PNN744,Q_PNN745,Q_PNN746,Q_PNN747,Q_PNN748,Q_PNN749,Q_PNN750,Q_PNN751,Q_PNN752,
             Q_PNN753,Q_PNN754,Q_PNN755;

wire PNN250,PNN251,PNN252,PNN253,PNN254,PNN255,PNN256,PNN257,PNN258,PNN259,
     PNN260,PNN261,PNN262,PNN263,PNN264,PNN265,PNN266,PNN267,PNN268,PNN269,
     PNN270,PNN271,PNN272,PNN273,PNN274,PNN275,PNN276,PNN277,PNN278,PNN279,
     PNN280,PNN281,PNN282,PNN283,PNN284,PNN285,PNN286,PNN287,PNN288,PNN289,
     PNN290,PNN293,PNN296,PNN299,PNN302,PNN305,PNN308,PNN311,PNN314,PNN315,
     PNN316,PNN317,PNN318,PNN319,PNN320,PNN321,PNN338,PNN339,PNN340,PNN341,
     PNN342,PNN343,PNN344,PNN345,PNN346,PNN347,PNN348,PNN349,PNN350,PNN351,
     PNN352,PNN353,PNN354,PNN367,PNN380,PNN393,PNN406,PNN419,PNN432,PNN445,
     PNN554,PNN555,PNN556,PNN557,PNN558,PNN559,PNN560,PNN561,PNN562,PNN563,
     PNN564,PNN565,PNN566,PNN567,PNN568,PNN569,PNN570,PNN571,PNN572,PNN573,
     PNN574,PNN575,PNN576,PNN577,PNN578,PNN579,PNN580,PNN581,PNN582,PNN583,
     PNN584,PNN585,PNN586,PNN587,PNN588,PNN589,PNN590,PNN591,PNN592,PNN593,
     PNN594,PNN595,PNN596,PNN597,PNN598,PNN599,PNN600,PNN601,PNN602,PNN607,
     PNN620,PNN625,PNN630,PNN635,PNN640,PNN645,PNN650,PNN655,PNN692,PNN693,
     PNN694,PNN695,PNN696,PNN697,PNN698,PNN699,PNN700,PNN701,PNN702,PNN703,
     PNN704,PNN705,PNN706,PNN707,PNN708,PNN709,PNN710,PNN711,PNN712,PNN713,
     PNN714,PNN715,PNN716,PNN717,PNN718,PNN719,PNN720,PNN721,PNN722,PNN723;

c499 c0 (IPNN_PNN1,IPNN_PNN5,IPNN_PNN9,IPNN_PNN13,IPNN_PNN17,IPNN_PNN21,IPNN_PNN25,IPNN_PNN29,IPNN_PNN33,IPNN_PNN37,
             IPNN_PNN41,IPNN_PNN45,IPNN_PNN49,IPNN_PNN53,IPNN_PNN57,IPNN_PNN61,IPNN_PNN65,IPNN_PNN69,IPNN_PNN73,IPNN_PNN77,
             IPNN_PNN81,IPNN_PNN85,IPNN_PNN89,IPNN_PNN93,IPNN_PNN97,IPNN_PNN101,IPNN_PNN105,IPNN_PNN109,IPNN_PNN113,IPNN_PNN117,
             IPNN_PNN121,IPNN_PNN125,IPNN_PNN129,IPNN_PNN130,IPNN_PNN131,IPNN_PNN132,IPNN_PNN133,IPNN_PNN134,IPNN_PNN135,IPNN_PNN136,
             IPNN_PNN137, PNN724,PNN725,PNN726,PNN727,PNN728,PNN729,PNN730,PNN731,PNN732,
             PNN733,PNN734,PNN735,PNN736,PNN737,PNN738,PNN739,PNN740,PNN741,PNN742,
             PNN743,PNN744,PNN745,PNN746,PNN747,PNN748,PNN749,PNN750,PNN751,PNN752,
             PNN753,PNN754,PNN755);


//Input FFs

dff iDFF_1  ( IPNN_PNN1  , PNN1, clk);
dff iDFF_2  ( IPNN_PNN5  , PNN5, clk);
dff iDFF_3  ( IPNN_PNN9  , PNN9, clk);
dff iDFF_4  ( IPNN_PNN13 , PNN13, clk);
dff iDFF_5  ( IPNN_PNN17 , PNN17, clk);
dff iDFF_6  ( IPNN_PNN21 , PNN21, clk);
dff iDFF_7  ( IPNN_PNN25 , PNN25, clk);
dff iDFF_8  ( IPNN_PNN29 , PNN29, clk);
dff iDFF_9  ( IPNN_PNN33 , PNN33, clk);
dff iDFF_10 ( IPNN_PNN37 , PNN37, clk);
dff iDFF_11 ( IPNN_PNN41 , PNN41, clk);
dff iDFF_12 ( IPNN_PNN45 , PNN45, clk);
dff iDFF_13 ( IPNN_PNN49 , PNN49, clk);
dff iDFF_14 ( IPNN_PNN53 , PNN53, clk);
dff iDFF_15 ( IPNN_PNN57 , PNN57, clk);
dff iDFF_16 ( IPNN_PNN61 , PNN61, clk);
dff iDFF_17 ( IPNN_PNN65 , PNN65, clk);
dff iDFF_18 ( IPNN_PNN69 , PNN69, clk);
dff iDFF_19 ( IPNN_PNN73 , PNN73, clk);
dff iDFF_20 ( IPNN_PNN77 , PNN77, clk);
dff iDFF_21 ( IPNN_PNN81 , PNN81, clk);
dff iDFF_22 ( IPNN_PNN85 , PNN85, clk);
dff iDFF_23 ( IPNN_PNN89 , PNN89, clk);
dff iDFF_24 ( IPNN_PNN93 , PNN93, clk);
dff iDFF_25 ( IPNN_PNN97 , PNN97, clk);
dff iDFF_26 ( IPNN_PNN101, PNN101, clk);
dff iDFF_27 ( IPNN_PNN105, PNN105, clk);
dff iDFF_28 ( IPNN_PNN109, PNN109, clk);
dff iDFF_29 ( IPNN_PNN113, PNN113, clk);
dff iDFF_30 ( IPNN_PNN117, PNN117, clk);
dff iDFF_31 ( IPNN_PNN121, PNN121, clk);
dff iDFF_32 ( IPNN_PNN125, PNN125, clk);
dff iDFF_33 ( IPNN_PNN129, PNN129, clk);
dff iDFF_34 ( IPNN_PNN130, PNN130, clk);
dff iDFF_35 ( IPNN_PNN131, PNN131, clk);
dff iDFF_36 ( IPNN_PNN132, PNN132, clk);
dff iDFF_37 ( IPNN_PNN133, PNN133, clk);
dff iDFF_38 ( IPNN_PNN134, PNN134, clk);
dff iDFF_39 ( IPNN_PNN135, PNN135, clk);
dff iDFF_40 ( IPNN_PNN136, PNN136, clk);
dff iDFF_41 ( IPNN_PNN137, PNN137, clk);


//output FFs
dff DFF_1 (Q_PNN724,PNN724,clk);
dff DFF_2 (Q_PNN725,PNN725,clk);
dff DFF_3 (Q_PNN726,PNN726,clk);
dff DFF_4 (Q_PNN727,PNN727,clk);
dff DFF_5 (Q_PNN728,PNN728,clk);
dff DFF_6 (Q_PNN729,PNN729,clk);
dff DFF_7 (Q_PNN730,PNN730,clk);
dff DFF_8 (Q_PNN731,PNN731,clk);
dff DFF_9 (Q_PNN732,PNN732,clk);
dff DFF_10(Q_PNN733,PNN733,clk);
dff DFF_11(Q_PNN734,PNN734,clk);
dff DFF_12(Q_PNN735,PNN735,clk);
dff DFF_13(Q_PNN736,PNN736,clk);
dff DFF_14(Q_PNN737,PNN737,clk);
dff DFF_15(Q_PNN738,PNN738,clk);
dff DFF_16(Q_PNN739,PNN739,clk);
dff DFF_17(Q_PNN740,PNN740,clk);
dff DFF_18(Q_PNN741,PNN741,clk);
dff DFF_19(Q_PNN742,PNN742,clk);
dff DFF_20(Q_PNN743,PNN743,clk);
dff DFF_21(Q_PNN744,PNN744,clk);
dff DFF_22(Q_PNN745,PNN745,clk);
dff DFF_23(Q_PNN746,PNN746,clk);
dff DFF_24(Q_PNN747,PNN747,clk);
dff DFF_25(Q_PNN748,PNN748,clk);
dff DFF_26(Q_PNN749,PNN749,clk);
dff DFF_27(Q_PNN750,PNN750,clk);
dff DFF_28(Q_PNN751,PNN751,clk);
dff DFF_29(Q_PNN752,PNN752,clk);
dff DFF_30(Q_PNN753,PNN753,clk);
dff DFF_31(Q_PNN754,PNN754,clk);
dff DFF_32(Q_PNN755,PNN755,clk);

endmodule
