
`timescale 1ns/100ps

module dff (q, d,clk);

input clk, d;
output q;
reg q;
always @(posedge clk) 
q = d;

endmodule


// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26

module c880 (PCN1,PCN8,PCN13,PCN17,PCN26,PCN29,PCN36,PCN42,PCN51,PCN55,
             PCN59,PCN68,PCN72,PCN73,PCN74,PCN75,PCN80,PCN85,PCN86,PCN87,
             PCN88,PCN89,PCN90,PCN91,PCN96,PCN101,PCN106,PCN111,PCN116,PCN121,
             PCN126,PCN130,PCN135,PCN138,PCN143,PCN146,PCN149,PCN152,PCN153,PCN156,
             PCN159,PCN165,PCN171,PCN177,PCN183,PCN189,PCN195,PCN201,PCN207,PCN210,
             PCN219,PCN228,PCN237,PCN246,PCN255,PCN259,PCN260,PCN261,PCN267,PCN268,
             PCN388,PCN389,PCN390,PCN391,PCN418,PCN419,PCN420,PCN421,PCN422,PCN423,
             PCN446,PCN447,PCN448,PCN449,PCN450,PCN767,PCN768,PCN850,PCN863,PCN864,
             PCN865,PCN866,PCN874,PCN878,PCN879,PCN880);

input PCN1,PCN8,PCN13,PCN17,PCN26,PCN29,PCN36,PCN42,PCN51,PCN55,
      PCN59,PCN68,PCN72,PCN73,PCN74,PCN75,PCN80,PCN85,PCN86,PCN87,
      PCN88,PCN89,PCN90,PCN91,PCN96,PCN101,PCN106,PCN111,PCN116,PCN121,
      PCN126,PCN130,PCN135,PCN138,PCN143,PCN146,PCN149,PCN152,PCN153,PCN156,
      PCN159,PCN165,PCN171,PCN177,PCN183,PCN189,PCN195,PCN201,PCN207,PCN210,
      PCN219,PCN228,PCN237,PCN246,PCN255,PCN259,PCN260,PCN261,PCN267,PCN268;

output PCN388,PCN389,PCN390,PCN391,PCN418,PCN419,PCN420,PCN421,PCN422,PCN423,
       PCN446,PCN447,PCN448,PCN449,PCN450,PCN767,PCN768,PCN850,PCN863,PCN864,
       PCN865,PCN866,PCN874,PCN878,PCN879,PCN880;

wire PCN269,PCN270,PCN273,PCN276,PCN279,PCN280,PCN284,PCN285,PCN286,PCN287,
     PCN290,PCN291,PCN292,PCN293,PCN294,PCN295,PCN296,PCN297,PCN298,PCN301,
     PCN302,PCN303,PCN304,PCN305,PCN306,PCN307,PCN308,PCN309,PCN310,PCN316,
     PCN317,PCN318,PCN319,PCN322,PCN323,PCN324,PCN325,PCN326,PCN327,PCN328,
     PCN329,PCN330,PCN331,PCN332,PCN333,PCN334,PCN335,PCN336,PCN337,PCN338,
     PCN339,PCN340,PCN341,PCN342,PCN343,PCN344,PCN345,PCN346,PCN347,PCN348,
     PCN349,PCN350,PCN351,PCN352,PCN353,PCN354,PCN355,PCN356,PCN357,PCN360,
     PCN363,PCN366,PCN369,PCN375,PCN376,PCN379,PCN382,PCN385,PCN392,PCN393,
     PCN399,PCN400,PCN401,PCN402,PCN403,PCN404,PCN405,PCN406,PCN407,PCN408,
     PCN409,PCN410,PCN411,PCN412,PCN413,PCN414,PCN415,PCN416,PCN417,PCN424,
     PCN425,PCN426,PCN427,PCN432,PCN437,PCN442,PCN443,PCN444,PCN445,PCN451,
     PCN460,PCN463,PCN466,PCN475,PCN476,PCN477,PCN478,PCN479,PCN480,PCN481,
     PCN482,PCN483,PCN488,PCN489,PCN490,PCN491,PCN492,PCN495,PCN498,PCN499,
     PCN500,PCN501,PCN502,PCN503,PCN504,PCN505,PCN506,PCN507,PCN508,PCN509,
     PCN510,PCN511,PCN512,PCN513,PCN514,PCN515,PCN516,PCN517,PCN518,PCN519,
     PCN520,PCN521,PCN522,PCN523,PCN524,PCN525,PCN526,PCN527,PCN528,PCN529,
     PCN530,PCN533,PCN536,PCN537,PCN538,PCN539,PCN540,PCN541,PCN542,PCN543,
     PCN544,PCN547,PCN550,PCN551,PCN552,PCN553,PCN557,PCN561,PCN565,PCN569,
     PCN573,PCN577,PCN581,PCN585,PCN586,PCN587,PCN588,PCN589,PCN590,PCN593,
     PCN596,PCN597,PCN600,PCN605,PCN606,PCN609,PCN615,PCN616,PCN619,PCN624,
     PCN625,PCN628,PCN631,PCN632,PCN635,PCN640,PCN641,PCN644,PCN650,PCN651,
     PCN654,PCN659,PCN660,PCN661,PCN662,PCN665,PCN669,PCN670,PCN673,PCN677,
     PCN678,PCN682,PCN686,PCN687,PCN692,PCN696,PCN697,PCN700,PCN704,PCN705,
     PCN708,PCN712,PCN713,PCN717,PCN721,PCN722,PCN727,PCN731,PCN732,PCN733,
     PCN734,PCN735,PCN736,PCN737,PCN738,PCN739,PCN740,PCN741,PCN742,PCN743,
     PCN744,PCN745,PCN746,PCN747,PCN748,PCN749,PCN750,PCN751,PCN752,PCN753,
     PCN754,PCN755,PCN756,PCN757,PCN758,PCN759,PCN760,PCN761,PCN762,PCN763,
     PCN764,PCN765,PCN766,PCN769,PCN770,PCN771,PCN772,PCN773,PCN777,PCN778,
     PCN781,PCN782,PCN785,PCN786,PCN787,PCN788,PCN789,PCN790,PCN791,PCN792,
     PCN793,PCN794,PCN795,PCN796,PCN802,PCN803,PCN804,PCN805,PCN806,PCN807,
     PCN808,PCN809,PCN810,PCN811,PCN812,PCN813,PCN814,PCN815,PCN819,PCN822,
     PCN825,PCN826,PCN827,PCN828,PCN829,PCN830,PCN831,PCN832,PCN833,PCN834,
     PCN835,PCN836,PCN837,PCN838,PCN839,PCN840,PCN841,PCN842,PCN843,PCN844,
     PCN845,PCN846,PCN847,PCN848,PCN849,PCN851,PCN852,PCN853,PCN854,PCN855,
     PCN856,PCN857,PCN858,PCN859,PCN860,PCN861,PCN862,PCN867,PCN868,PCN869,
     PCN870,PCN871,PCN872,PCN873,PCN875,PCN876,PCN877;

nand NAND4_1 (PCN269, PCN1, PCN8, PCN13, PCN17);
nand NAND4_2 (PCN270, PCN1, PCN26, PCN13, PCN17);
and AND3_3 (PCN273, PCN29, PCN36, PCN42);
and AND3_4 (PCN276, PCN1, PCN26, PCN51);
nand NAND4_5 (PCN279, PCN1, PCN8, PCN51, PCN17);
nand NAND4_6 (PCN280, PCN1, PCN8, PCN13, PCN55);
nand NAND4_7 (PCN284, PCN59, PCN42, PCN68, PCN72);
nand NAND2_8 (PCN285, PCN29, PCN68);
nand NAND3_9 (PCN286, PCN59, PCN68, PCN74);
and AND3_10 (PCN287, PCN29, PCN75, PCN80);
and AND3_11 (PCN290, PCN29, PCN75, PCN42);
and AND3_12 (PCN291, PCN29, PCN36, PCN80);
and AND3_13 (PCN292, PCN29, PCN36, PCN42);
and AND3_14 (PCN293, PCN59, PCN75, PCN80);
and AND3_15 (PCN294, PCN59, PCN75, PCN42);
and AND3_16 (PCN295, PCN59, PCN36, PCN80);
and AND3_17 (PCN296, PCN59, PCN36, PCN42);
and AND2_18 (PCN297, PCN85, PCN86);
or OR2_19 (PCN298, PCN87, PCN88);
nand NAND2_20 (PCN301, PCN91, PCN96);
or OR2_21 (PCN302, PCN91, PCN96);
nand NAND2_22 (PCN303, PCN101, PCN106);
or OR2_23 (PCN304, PCN101, PCN106);
nand NAND2_24 (PCN305, PCN111, PCN116);
or OR2_25 (PCN306, PCN111, PCN116);
nand NAND2_26 (PCN307, PCN121, PCN126);
or OR2_27 (PCN308, PCN121, PCN126);
and AND2_28 (PCN309, PCN8, PCN138);
not NOT1_29 (PCN310, PCN268);
and AND2_30 (PCN316, PCN51, PCN138);
and AND2_31 (PCN317, PCN17, PCN138);
and AND2_32 (PCN318, PCN152, PCN138);
nand NAND2_33 (PCN319, PCN59, PCN156);
nor NOR2_34 (PCN322, PCN17, PCN42);
and AND2_35 (PCN323, PCN17, PCN42);
nand NAND2_36 (PCN324, PCN159, PCN165);
or OR2_37 (PCN325, PCN159, PCN165);
nand NAND2_38 (PCN326, PCN171, PCN177);
or OR2_39 (PCN327, PCN171, PCN177);
nand NAND2_40 (PCN328, PCN183, PCN189);
or OR2_41 (PCN329, PCN183, PCN189);
nand NAND2_42 (PCN330, PCN195, PCN201);
or OR2_43 (PCN331, PCN195, PCN201);
and AND2_44 (PCN332, PCN210, PCN91);
and AND2_45 (PCN333, PCN210, PCN96);
and AND2_46 (PCN334, PCN210, PCN101);
and AND2_47 (PCN335, PCN210, PCN106);
and AND2_48 (PCN336, PCN210, PCN111);
and AND2_49 (PCN337, PCN255, PCN259);
and AND2_50 (PCN338, PCN210, PCN116);
and AND2_51 (PCN339, PCN255, PCN260);
and AND2_52 (PCN340, PCN210, PCN121);
and AND2_53 (PCN341, PCN255, PCN267);
not NOT1_54 (PCN342, PCN269);
not NOT1_55 (PCN343, PCN273);
or OR2_56 (PCN344, PCN270, PCN273);
not NOT1_57 (PCN345, PCN276);
not NOT1_58 (PCN346, PCN276);
not NOT1_59 (PCN347, PCN279);
nor NOR2_60 (PCN348, PCN280, PCN284);
or OR2_61 (PCN349, PCN280, PCN285);
or OR2_62 (PCN350, PCN280, PCN286);
not NOT1_63 (PCN351, PCN293);
not NOT1_64 (PCN352, PCN294);
not NOT1_65 (PCN353, PCN295);
not NOT1_66 (PCN354, PCN296);
nand NAND2_67 (PCN355, PCN89, PCN298);
and AND2_68 (PCN356, PCN90, PCN298);
nand NAND2_69 (PCN357, PCN301, PCN302);
nand NAND2_70 (PCN360, PCN303, PCN304);
nand NAND2_71 (PCN363, PCN305, PCN306);
nand NAND2_72 (PCN366, PCN307, PCN308);
not NOT1_73 (PCN369, PCN310);
nor NOR2_74 (PCN375, PCN322, PCN323);
nand NAND2_75 (PCN376, PCN324, PCN325);
nand NAND2_76 (PCN379, PCN326, PCN327);
nand NAND2_77 (PCN382, PCN328, PCN329);
nand NAND2_78 (PCN385, PCN330, PCN331);
buf BUFF1_79 (PCN388, PCN290);
buf BUFF1_80 (PCN389, PCN291);
buf BUFF1_81 (PCN390, PCN292);
buf BUFF1_82 (PCN391, PCN297);
or OR2_83 (PCN392, PCN270, PCN343);
not NOT1_84 (PCN393, PCN345);
not NOT1_85 (PCN399, PCN346);
and AND2_86 (PCN400, PCN348, PCN73);
not NOT1_87 (PCN401, PCN349);
not NOT1_88 (PCN402, PCN350);
not NOT1_89 (PCN403, PCN355);
not NOT1_90 (PCN404, PCN357);
not NOT1_91 (PCN405, PCN360);
and AND2_92 (PCN406, PCN357, PCN360);
not NOT1_93 (PCN407, PCN363);
not NOT1_94 (PCN408, PCN366);
and AND2_95 (PCN409, PCN363, PCN366);
nand NAND2_96 (PCN410, PCN347, PCN352);
not NOT1_97 (PCN411, PCN376);
not NOT1_98 (PCN412, PCN379);
and AND2_99 (PCN413, PCN376, PCN379);
not NOT1_100 (PCN414, PCN382);
not NOT1_101 (PCN415, PCN385);
and AND2_102 (PCN416, PCN382, PCN385);
and AND2_103 (PCN417, PCN210, PCN369);
buf BUFF1_104 (PCN418, PCN342);
buf BUFF1_105 (PCN419, PCN344);
buf BUFF1_106 (PCN420, PCN351);
buf BUFF1_107 (PCN421, PCN353);
buf BUFF1_108 (PCN422, PCN354);
buf BUFF1_109 (PCN423, PCN356);
not NOT1_110 (PCN424, PCN400);
and AND2_111 (PCN425, PCN404, PCN405);
and AND2_112 (PCN426, PCN407, PCN408);
and AND3_113 (PCN427, PCN319, PCN393, PCN55);
and AND3_114 (PCN432, PCN393, PCN17, PCN287);
nand NAND3_115 (PCN437, PCN393, PCN287, PCN55);
nand NAND4_116 (PCN442, PCN375, PCN59, PCN156, PCN393);
nand NAND3_117 (PCN443, PCN393, PCN319, PCN17);
and AND2_118 (PCN444, PCN411, PCN412);
and AND2_119 (PCN445, PCN414, PCN415);
buf BUFF1_120 (PCN446, PCN392);
buf BUFF1_121 (PCN447, PCN399);
buf BUFF1_122 (PCN448, PCN401);
buf BUFF1_123 (PCN449, PCN402);
buf BUFF1_124 (PCN450, PCN403);
not NOT1_125 (PCN451, PCN424);
nor NOR2_126 (PCN460, PCN406, PCN425);
nor NOR2_127 (PCN463, PCN409, PCN426);
nand NAND2_128 (PCN466, PCN442, PCN410);
and AND2_129 (PCN475, PCN143, PCN427);
and AND2_130 (PCN476, PCN310, PCN432);
and AND2_131 (PCN477, PCN146, PCN427);
and AND2_132 (PCN478, PCN310, PCN432);
and AND2_133 (PCN479, PCN149, PCN427);
and AND2_134 (PCN480, PCN310, PCN432);
and AND2_135 (PCN481, PCN153, PCN427);
and AND2_136 (PCN482, PCN310, PCN432);
nand NAND2_137 (PCN483, PCN443, PCN1);
or OR2_138 (PCN488, PCN369, PCN437);
or OR2_139 (PCN489, PCN369, PCN437);
or OR2_140 (PCN490, PCN369, PCN437);
or OR2_141 (PCN491, PCN369, PCN437);
nor NOR2_142 (PCN492, PCN413, PCN444);
nor NOR2_143 (PCN495, PCN416, PCN445);
nand NAND2_144 (PCN498, PCN130, PCN460);
or OR2_145 (PCN499, PCN130, PCN460);
nand NAND2_146 (PCN500, PCN463, PCN135);
or OR2_147 (PCN501, PCN463, PCN135);
and AND2_148 (PCN502, PCN91, PCN466);
nor NOR2_149 (PCN503, PCN475, PCN476);
and AND2_150 (PCN504, PCN96, PCN466);
nor NOR2_151 (PCN505, PCN477, PCN478);
and AND2_152 (PCN506, PCN101, PCN466);
nor NOR2_153 (PCN507, PCN479, PCN480);
and AND2_154 (PCN508, PCN106, PCN466);
nor NOR2_155 (PCN509, PCN481, PCN482);
and AND2_156 (PCN510, PCN143, PCN483);
and AND2_157 (PCN511, PCN111, PCN466);
and AND2_158 (PCN512, PCN146, PCN483);
and AND2_159 (PCN513, PCN116, PCN466);
and AND2_160 (PCN514, PCN149, PCN483);
and AND2_161 (PCN515, PCN121, PCN466);
and AND2_162 (PCN516, PCN153, PCN483);
and AND2_163 (PCN517, PCN126, PCN466);
nand NAND2_164 (PCN518, PCN130, PCN492);
or OR2_165 (PCN519, PCN130, PCN492);
nand NAND2_166 (PCN520, PCN495, PCN207);
or OR2_167 (PCN521, PCN495, PCN207);
and AND2_168 (PCN522, PCN451, PCN159);
and AND2_169 (PCN523, PCN451, PCN165);
and AND2_170 (PCN524, PCN451, PCN171);
and AND2_171 (PCN525, PCN451, PCN177);
and AND2_172 (PCN526, PCN451, PCN183);
nand NAND2_173 (PCN527, PCN451, PCN189);
nand NAND2_174 (PCN528, PCN451, PCN195);
nand NAND2_175 (PCN529, PCN451, PCN201);
nand NAND2_176 (PCN530, PCN498, PCN499);
nand NAND2_177 (PCN533, PCN500, PCN501);
nor NOR2_178 (PCN536, PCN309, PCN502);
nor NOR2_179 (PCN537, PCN316, PCN504);
nor NOR2_180 (PCN538, PCN317, PCN506);
nor NOR2_181 (PCN539, PCN318, PCN508);
nor NOR2_182 (PCN540, PCN510, PCN511);
nor NOR2_183 (PCN541, PCN512, PCN513);
nor NOR2_184 (PCN542, PCN514, PCN515);
nor NOR2_185 (PCN543, PCN516, PCN517);
nand NAND2_186 (PCN544, PCN518, PCN519);
nand NAND2_187 (PCN547, PCN520, PCN521);
not NOT1_188 (PCN550, PCN530);
not NOT1_189 (PCN551, PCN533);
and AND2_190 (PCN552, PCN530, PCN533);
nand NAND2_191 (PCN553, PCN536, PCN503);
nand NAND2_192 (PCN557, PCN537, PCN505);
nand NAND2_193 (PCN561, PCN538, PCN507);
nand NAND2_194 (PCN565, PCN539, PCN509);
nand NAND2_195 (PCN569, PCN488, PCN540);
nand NAND2_196 (PCN573, PCN489, PCN541);
nand NAND2_197 (PCN577, PCN490, PCN542);
nand NAND2_198 (PCN581, PCN491, PCN543);
not NOT1_199 (PCN585, PCN544);
not NOT1_200 (PCN586, PCN547);
and AND2_201 (PCN587, PCN544, PCN547);
and AND2_202 (PCN588, PCN550, PCN551);
and AND2_203 (PCN589, PCN585, PCN586);
nand NAND2_204 (PCN590, PCN553, PCN159);
or OR2_205 (PCN593, PCN553, PCN159);
and AND2_206 (PCN596, PCN246, PCN553);
nand NAND2_207 (PCN597, PCN557, PCN165);
or OR2_208 (PCN600, PCN557, PCN165);
and AND2_209 (PCN605, PCN246, PCN557);
nand NAND2_210 (PCN606, PCN561, PCN171);
or OR2_211 (PCN609, PCN561, PCN171);
and AND2_212 (PCN615, PCN246, PCN561);
nand NAND2_213 (PCN616, PCN565, PCN177);
or OR2_214 (PCN619, PCN565, PCN177);
and AND2_215 (PCN624, PCN246, PCN565);
nand NAND2_216 (PCN625, PCN569, PCN183);
or OR2_217 (PCN628, PCN569, PCN183);
and AND2_218 (PCN631, PCN246, PCN569);
nand NAND2_219 (PCN632, PCN573, PCN189);
or OR2_220 (PCN635, PCN573, PCN189);
and AND2_221 (PCN640, PCN246, PCN573);
nand NAND2_222 (PCN641, PCN577, PCN195);
or OR2_223 (PCN644, PCN577, PCN195);
and AND2_224 (PCN650, PCN246, PCN577);
nand NAND2_225 (PCN651, PCN581, PCN201);
or OR2_226 (PCN654, PCN581, PCN201);
and AND2_227 (PCN659, PCN246, PCN581);
nor NOR2_228 (PCN660, PCN552, PCN588);
nor NOR2_229 (PCN661, PCN587, PCN589);
not NOT1_230 (PCN662, PCN590);
and AND2_231 (PCN665, PCN593, PCN590);
nor NOR2_232 (PCN669, PCN596, PCN522);
not NOT1_233 (PCN670, PCN597);
and AND2_234 (PCN673, PCN600, PCN597);
nor NOR2_235 (PCN677, PCN605, PCN523);
not NOT1_236 (PCN678, PCN606);
and AND2_237 (PCN682, PCN609, PCN606);
nor NOR2_238 (PCN686, PCN615, PCN524);
not NOT1_239 (PCN687, PCN616);
and AND2_240 (PCN692, PCN619, PCN616);
nor NOR2_241 (PCN696, PCN624, PCN525);
not NOT1_242 (PCN697, PCN625);
and AND2_243 (PCN700, PCN628, PCN625);
nor NOR2_244 (PCN704, PCN631, PCN526);
not NOT1_245 (PCN705, PCN632);
and AND2_246 (PCN708, PCN635, PCN632);
nor NOR2_247 (PCN712, PCN337, PCN640);
not NOT1_248 (PCN713, PCN641);
and AND2_249 (PCN717, PCN644, PCN641);
nor NOR2_250 (PCN721, PCN339, PCN650);
not NOT1_251 (PCN722, PCN651);
and AND2_252 (PCN727, PCN654, PCN651);
nor NOR2_253 (PCN731, PCN341, PCN659);
nand NAND2_254 (PCN732, PCN654, PCN261);
nand NAND3_255 (PCN733, PCN644, PCN654, PCN261);
nand NAND4_256 (PCN734, PCN635, PCN644, PCN654, PCN261);
not NOT1_257 (PCN735, PCN662);
and AND2_258 (PCN736, PCN228, PCN665);
and AND2_259 (PCN737, PCN237, PCN662);
not NOT1_260 (PCN738, PCN670);
and AND2_261 (PCN739, PCN228, PCN673);
and AND2_262 (PCN740, PCN237, PCN670);
not NOT1_263 (PCN741, PCN678);
and AND2_264 (PCN742, PCN228, PCN682);
and AND2_265 (PCN743, PCN237, PCN678);
not NOT1_266 (PCN744, PCN687);
and AND2_267 (PCN745, PCN228, PCN692);
and AND2_268 (PCN746, PCN237, PCN687);
not NOT1_269 (PCN747, PCN697);
and AND2_270 (PCN748, PCN228, PCN700);
and AND2_271 (PCN749, PCN237, PCN697);
not NOT1_272 (PCN750, PCN705);
and AND2_273 (PCN751, PCN228, PCN708);
and AND2_274 (PCN752, PCN237, PCN705);
not NOT1_275 (PCN753, PCN713);
and AND2_276 (PCN754, PCN228, PCN717);
and AND2_277 (PCN755, PCN237, PCN713);
not NOT1_278 (PCN756, PCN722);
nor NOR2_279 (PCN757, PCN727, PCN261);
and AND2_280 (PCN758, PCN727, PCN261);
and AND2_281 (PCN759, PCN228, PCN727);
and AND2_282 (PCN760, PCN237, PCN722);
nand NAND2_283 (PCN761, PCN644, PCN722);
nand NAND2_284 (PCN762, PCN635, PCN713);
nand NAND3_285 (PCN763, PCN635, PCN644, PCN722);
nand NAND2_286 (PCN764, PCN609, PCN687);
nand NAND2_287 (PCN765, PCN600, PCN678);
nand NAND3_288 (PCN766, PCN600, PCN609, PCN687);
buf BUFF1_289 (PCN767, PCN660);
buf BUFF1_290 (PCN768, PCN661);
nor NOR2_291 (PCN769, PCN736, PCN737);
nor NOR2_292 (PCN770, PCN739, PCN740);
nor NOR2_293 (PCN771, PCN742, PCN743);
nor NOR2_294 (PCN772, PCN745, PCN746);
nand NAND4_295 (PCN773, PCN750, PCN762, PCN763, PCN734);
nor NOR2_296 (PCN777, PCN748, PCN749);
nand NAND3_297 (PCN778, PCN753, PCN761, PCN733);
nor NOR2_298 (PCN781, PCN751, PCN752);
nand NAND2_299 (PCN782, PCN756, PCN732);
nor NOR2_300 (PCN785, PCN754, PCN755);
nor NOR2_301 (PCN786, PCN757, PCN758);
nor NOR2_302 (PCN787, PCN759, PCN760);
nor NOR2_303 (PCN788, PCN700, PCN773);
and AND2_304 (PCN789, PCN700, PCN773);
nor NOR2_305 (PCN790, PCN708, PCN778);
and AND2_306 (PCN791, PCN708, PCN778);
nor NOR2_307 (PCN792, PCN717, PCN782);
and AND2_308 (PCN793, PCN717, PCN782);
and AND2_309 (PCN794, PCN219, PCN786);
nand NAND2_310 (PCN795, PCN628, PCN773);
nand NAND2_311 (PCN796, PCN795, PCN747);
nor NOR2_312 (PCN802, PCN788, PCN789);
nor NOR2_313 (PCN803, PCN790, PCN791);
nor NOR2_314 (PCN804, PCN792, PCN793);
nor NOR2_315 (PCN805, PCN340, PCN794);
nor NOR2_316 (PCN806, PCN692, PCN796);
and AND2_317 (PCN807, PCN692, PCN796);
and AND2_318 (PCN808, PCN219, PCN802);
and AND2_319 (PCN809, PCN219, PCN803);
and AND2_320 (PCN810, PCN219, PCN804);
nand NAND4_321 (PCN811, PCN805, PCN787, PCN731, PCN529);
nand NAND2_322 (PCN812, PCN619, PCN796);
nand NAND3_323 (PCN813, PCN609, PCN619, PCN796);
nand NAND4_324 (PCN814, PCN600, PCN609, PCN619, PCN796);
nand NAND4_325 (PCN815, PCN738, PCN765, PCN766, PCN814);
nand NAND3_326 (PCN819, PCN741, PCN764, PCN813);
nand NAND2_327 (PCN822, PCN744, PCN812);
nor NOR2_328 (PCN825, PCN806, PCN807);
nor NOR2_329 (PCN826, PCN335, PCN808);
nor NOR2_330 (PCN827, PCN336, PCN809);
nor NOR2_331 (PCN828, PCN338, PCN810);
not NOT1_332 (PCN829, PCN811);
nor NOR2_333 (PCN830, PCN665, PCN815);
and AND2_334 (PCN831, PCN665, PCN815);
nor NOR2_335 (PCN832, PCN673, PCN819);
and AND2_336 (PCN833, PCN673, PCN819);
nor NOR2_337 (PCN834, PCN682, PCN822);
and AND2_338 (PCN835, PCN682, PCN822);
and AND2_339 (PCN836, PCN219, PCN825);
nand NAND3_340 (PCN837, PCN826, PCN777, PCN704);
nand NAND4_341 (PCN838, PCN827, PCN781, PCN712, PCN527);
nand NAND4_342 (PCN839, PCN828, PCN785, PCN721, PCN528);
not NOT1_343 (PCN840, PCN829);
nand NAND2_344 (PCN841, PCN815, PCN593);
nor NOR2_345 (PCN842, PCN830, PCN831);
nor NOR2_346 (PCN843, PCN832, PCN833);
nor NOR2_347 (PCN844, PCN834, PCN835);
nor NOR2_348 (PCN845, PCN334, PCN836);
not NOT1_349 (PCN846, PCN837);
not NOT1_350 (PCN847, PCN838);
not NOT1_351 (PCN848, PCN839);
and AND2_352 (PCN849, PCN735, PCN841);
buf BUFF1_353 (PCN850, PCN840);
and AND2_354 (PCN851, PCN219, PCN842);
and AND2_355 (PCN852, PCN219, PCN843);
and AND2_356 (PCN853, PCN219, PCN844);
nand NAND3_357 (PCN854, PCN845, PCN772, PCN696);
not NOT1_358 (PCN855, PCN846);
not NOT1_359 (PCN856, PCN847);
not NOT1_360 (PCN857, PCN848);
not NOT1_361 (PCN858, PCN849);
nor NOR2_362 (PCN859, PCN417, PCN851);
nor NOR2_363 (PCN860, PCN332, PCN852);
nor NOR2_364 (PCN861, PCN333, PCN853);
not NOT1_365 (PCN862, PCN854);
buf BUFF1_366 (PCN863, PCN855);
buf BUFF1_367 (PCN864, PCN856);
buf BUFF1_368 (PCN865, PCN857);
buf BUFF1_369 (PCN866, PCN858);
nand NAND3_370 (PCN867, PCN859, PCN769, PCN669);
nand NAND3_371 (PCN868, PCN860, PCN770, PCN677);
nand NAND3_372 (PCN869, PCN861, PCN771, PCN686);
not NOT1_373 (PCN870, PCN862);
not NOT1_374 (PCN871, PCN867);
not NOT1_375 (PCN872, PCN868);
not NOT1_376 (PCN873, PCN869);
buf BUFF1_377 (PCN874, PCN870);
not NOT1_378 (PCN875, PCN871);
not NOT1_379 (PCN876, PCN872);
not NOT1_380 (PCN877, PCN873);
buf BUFF1_381 (PCN878, PCN875);
buf BUFF1_382 (PCN879, PCN876);
buf BUFF1_383 (PCN880, PCN877);

endmodule



module c880_clk_ipFF (clk,PCN1,PCN8,PCN13,PCN17,PCN26,PCN29,PCN36,PCN42,PCN51,PCN55,
             PCN59,PCN68,PCN72,PCN73,PCN74,PCN75,PCN80,PCN85,PCN86,PCN87,
             PCN88,PCN89,PCN90,PCN91,PCN96,PCN101,PCN106,PCN111,PCN116,PCN121,
             PCN126,PCN130,PCN135,PCN138,PCN143,PCN146,PCN149,PCN152,PCN153,PCN156,
             PCN159,PCN165,PCN171,PCN177,PCN183,PCN189,PCN195,PCN201,PCN207,PCN210,
             PCN219,PCN228,PCN237,PCN246,PCN255,PCN259,PCN260,PCN261,PCN267,PCN268,
             Q_PCN388,Q_PCN389,Q_PCN390,Q_PCN391,Q_PCN418,Q_PCN419,Q_PCN420,Q_PCN421,Q_PCN422,Q_PCN423,
             Q_PCN446,Q_PCN447,Q_PCN448,Q_PCN449,Q_PCN450,Q_PCN767,Q_PCN768,Q_PCN850,Q_PCN863,Q_PCN864,
             Q_PCN865,Q_PCN866,Q_PCN874,Q_PCN878,Q_PCN879,Q_PCN880);

input clk,PCN1,PCN8,PCN13,PCN17,PCN26,PCN29,PCN36,PCN42,PCN51,PCN55,
      PCN59,PCN68,PCN72,PCN73,PCN74,PCN75,PCN80,PCN85,PCN86,PCN87,
      PCN88,PCN89,PCN90,PCN91,PCN96,PCN101,PCN106,PCN111,PCN116,PCN121,
      PCN126,PCN130,PCN135,PCN138,PCN143,PCN146,PCN149,PCN152,PCN153,PCN156,
      PCN159,PCN165,PCN171,PCN177,PCN183,PCN189,PCN195,PCN201,PCN207,PCN210,
      PCN219,PCN228,PCN237,PCN246,PCN255,PCN259,PCN260,PCN261,PCN267,PCN268;

output  Q_PCN388,Q_PCN389,Q_PCN390,Q_PCN391,Q_PCN418,Q_PCN419,Q_PCN420,Q_PCN421,Q_PCN422,Q_PCN423,
             Q_PCN446,Q_PCN447,Q_PCN448,Q_PCN449,Q_PCN450,Q_PCN767,Q_PCN768,Q_PCN850,Q_PCN863,Q_PCN864,
             Q_PCN865,Q_PCN866,Q_PCN874,Q_PCN878,Q_PCN879,Q_PCN880;

c880 c1 (INP_PCN1,INP_PCN8,INP_PCN13,INP_PCN17,INP_PCN26,INP_PCN29,INP_PCN36,INP_PCN42,INP_PCN51,INP_PCN55,
             INP_PCN59,INP_PCN68,INP_PCN72,INP_PCN73,INP_PCN74,INP_PCN75,INP_PCN80,INP_PCN85,INP_PCN86,INP_PCN87,
             INP_PCN88,INP_PCN89,INP_PCN90,INP_PCN91,INP_PCN96,INP_PCN101,INP_PCN106,INP_PCN111,INP_PCN116,INP_PCN121,
             INP_PCN126,INP_PCN130,INP_PCN135,INP_PCN138,INP_PCN143,INP_PCN146,INP_PCN149,INP_PCN152,INP_PCN153,INP_PCN156,
             INP_PCN159,INP_PCN165,INP_PCN171,INP_PCN177,INP_PCN183,INP_PCN189,INP_PCN195,INP_PCN201,INP_PCN207,INP_PCN210,
             INP_PCN219,INP_PCN228,INP_PCN237,INP_PCN246,INP_PCN255,INP_PCN259,INP_PCN260,INP_PCN261,INP_PCN267,INP_PCN268,          
             PCN388,PCN389,PCN390,PCN391,PCN418,PCN419,PCN420,PCN421,PCN422,PCN423,
             PCN446,PCN447,PCN448,PCN449,PCN450,PCN767,PCN768,PCN850,PCN863,PCN864,
             PCN865,PCN866,PCN874,PCN878,PCN879,PCN880);

//Input FFs
dff iDFF_1( INP_PCN1,  PCN1, clk);
dff iDFF_2( INP_PCN8,  PCN8, clk);
dff iDFF_3( INP_PCN13, PCN13,clk);
dff iDFF_4( INP_PCN17, PCN17,clk);
dff iDFF_5( INP_PCN26, PCN26,clk);
dff iDFF_6( INP_PCN29, PCN29,clk);
dff iDFF_7( INP_PCN36, PCN36,clk);
dff iDFF_8( INP_PCN42, PCN42,clk);
dff iDFF_9( INP_PCN51, PCN51,clk);
dff iDFF_10( INP_PCN55, PCN55,clk);
dff iDFF_11( INP_PCN59, PCN59,clk);
dff iDFF_12( INP_PCN68, PCN68,clk);
dff iDFF_13( INP_PCN72, PCN72,clk);
dff iDFF_14( INP_PCN73, PCN73,clk);
dff iDFF_15( INP_PCN74, PCN74,clk);
dff iDFF_16( INP_PCN75, PCN75,clk);
dff iDFF_17( INP_PCN80, PCN80,clk);
dff iDFF_18( INP_PCN85, PCN85,clk);
dff iDFF_19( INP_PCN86, PCN86,clk);
dff iDFF_20( INP_PCN87, PCN87,clk);
dff iDFF_21( INP_PCN88, PCN88,clk);
dff iDFF_22( INP_PCN89, PCN89,clk);
dff iDFF_23( INP_PCN90, PCN90,clk);
dff iDFF_24( INP_PCN91, PCN91,clk);
dff iDFF_25( INP_PCN96, PCN96,clk);
dff iDFF_26( INP_PCN101,PCN101,clk);
dff iDFF_27( INP_PCN106,PCN106,clk);
dff iDFF_28( INP_PCN111,PCN111,clk);
dff iDFF_29( INP_PCN116,PCN116,clk);
dff iDFF_30( INP_PCN121,PCN121,clk);
dff iDFF_31( INP_PCN126,PCN126,clk);
dff iDFF_32( INP_PCN130,PCN130,clk);
dff iDFF_33( INP_PCN135,PCN135,clk);
dff iDFF_34( INP_PCN138,PCN138,clk);
dff iDFF_35( INP_PCN143,PCN143,clk);
dff iDFF_36( INP_PCN146,PCN146,clk);
dff iDFF_37( INP_PCN149,PCN149,clk);
dff iDFF_38( INP_PCN152,PCN152,clk);
dff iDFF_39( INP_PCN153,PCN153,clk);
dff iDFF_40( INP_PCN156,PCN156,clk);
dff iDFF_41( INP_PCN159,PCN159,clk);
dff iDFF_42( INP_PCN165,PCN165,clk);
dff iDFF_43( INP_PCN171,PCN171,clk);
dff iDFF_44( INP_PCN177,PCN177,clk);
dff iDFF_45( INP_PCN183,PCN183,clk);
dff iDFF_46( INP_PCN189,PCN189,clk);
dff iDFF_47( INP_PCN195,PCN195,clk);
dff iDFF_48( INP_PCN201,PCN201,clk);
dff iDFF_49( INP_PCN207,PCN207,clk);
dff iDFF_50( INP_PCN210,PCN210,clk);
dff iDFF_51( INP_PCN219,PCN219,clk);
dff iDFF_52( INP_PCN228,PCN228,clk);
dff iDFF_53( INP_PCN237,PCN237,clk);
dff iDFF_54( INP_PCN246,PCN246,clk);
dff iDFF_55( INP_PCN255,PCN255,clk);
dff iDFF_56( INP_PCN259,PCN259,clk);
dff iDFF_57( INP_PCN260,PCN260,clk);
dff iDFF_58( INP_PCN261,PCN261,clk);
dff iDFF_59( INP_PCN267,PCN267,clk);
dff iDFF_60( INP_PCN268,PCN268,clk);

//Output FFs
dff DFF_1 (Q_PCN388,PCN388,clk);
dff DFF_2 (Q_PCN389,PCN389,clk);
dff DFF_3 (Q_PCN390,PCN390,clk);
dff DFF_4 (Q_PCN391,PCN391,clk);
dff DFF_5 (Q_PCN418,PCN418,clk);
dff DFF_6 (Q_PCN419,PCN419,clk);
dff DFF_7 (Q_PCN420,PCN420,clk);
dff DFF_8 (Q_PCN421,PCN421,clk);
dff DFF_9 (Q_PCN422,PCN422,clk);
dff DFF_10(Q_PCN423,PCN423,clk);
dff DFF_11(Q_PCN446,PCN446,clk);
dff DFF_12(Q_PCN447,PCN447,clk);
dff DFF_13(Q_PCN448,PCN448,clk);
dff DFF_14(Q_PCN449,PCN449,clk);
dff DFF_15(Q_PCN450,PCN450,clk);
dff DFF_16(Q_PCN767,PCN767,clk);
dff DFF_17(Q_PCN768,PCN768,clk);
dff DFF_18(Q_PCN850,PCN850,clk);
dff DFF_19(Q_PCN863,PCN863,clk);
dff DFF_20(Q_PCN864,PCN864,clk);
dff DFF_22(Q_PCN865,PCN865,clk);
dff DFF_23(Q_PCN866,PCN866,clk);
dff DFF_24(Q_PCN874,PCN874,clk);
dff DFF_25(Q_PCN878,PCN878,clk);
dff DFF_26(Q_PCN879,PCN879,clk);
dff DFF_27(Q_PCN880, PCN880,clk);


endmodule
