
.SUBCKT HS65_GSS1_FA1X21 A0 B0 CI CO S0 gnd gnds vdd vdds
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070516.0 at 17:38 5 Jun 2007
Xld_D0 gnds:F20 vdds:F21 DNWPS AREA=7.83275 PJ=13.5
MMM11 na:F43 A0:F44 gnd:F45 gnds:F42 NSVTGP W=0.67u L=0.06u 
MMM18 na:F103 A0:F104 vdd:F105 vdds:F102 PSVTGP W=1.02u L=0.06u 
MMM24 axorb:F29 na:F28 B0:F27 gnds:F26 NSVTGP W=0.48u L=0.06u 
MMM25 axorb:F89 A0:F88 B0:F87 vdds:F86 PSVTGP W=0.77u L=0.06u 
MMM28 axorb:F83 na:F84 nb:F85 vdds:F82 PSVTGP W=0.77u L=0.06u 
MMM29 axorb:F23 A0:F24 nb:F25 gnds:F22 NSVTGP W=0.48u L=0.06u 
MMM30 axnorb:F37 na:F36 nb:F35 gnds:F34 NSVTGP W=0.48u L=0.06u 
MMM31 axnorb:F97 A0:F96 nb:F95 vdds:F94 PSVTGP W=0.67u L=0.06u 
MMM32 axnorb:F91 na:F92 B0:F93 vdds:F90 PSVTGP W=0.89u L=0.06u 
MMM33 axnorb:F31 A0:F32 B0:F33 gnds:F30 NSVTGP W=0.43u L=0.06u 
MMM34 s:F55 axnorb:F56 net199:F57 gnds:F54 NSVTGP W=0.46u L=0.06u 
MMM35 s:F115 axorb:F116 net199:F117 vdds:F114 PSVTGP W=0.67u L=0.06u 
MMM36 s:F121 axnorb:F120 CI:F119 vdds:F118 PSVTGP W=0.81u L=0.06u 
MMM37 s:F61 axorb:F60 CI:F59 gnds:F58 NSVTGP W=0.47u L=0.06u 
MMM38 co1:F53 axorb:F52 net199:F51 gnds:F50 NSVTGP W=0.46u L=0.06u 
MMM39 co1:F113 axnorb:F112 net199:F111 vdds:F110 PSVTGP W=0.51u L=0.06u 
MMM40 co1:F107 axorb:F108 na:F109 vdds:F106 PSVTGP W=0.51u L=0.06u 
MMM41 co1:F47 axnorb:F48 na:F49 gnds:F46 NSVTGP W=0.46u L=0.06u 
MMM50 nb:F41 B0:F40 gnd:F39 gnds:F38 NSVTGP W=0.48u L=0.06u 
MMM51 nb:F101 B0:F100 vdd:F99 vdds:F98 PSVTGP W=0.67u L=0.06u 
MMM52 net199:F65 CI:F64 gnd:F63 gnds:F62 NSVTGP W=0.46u L=0.06u 
MMM53 net199:F125 CI:F124 vdd:F123 vdds:F122 PSVTGP W=0.74u L=0.06u 
MMM56 S0:F67 s:F68 gnd:F69 gnds:F66 NSVTGP W=0.77u L=0.06u 
MMM56@2 S0:F73 s:F72 gnd:F71 gnds:F70 NSVTGP W=0.77u L=0.06u 
MMM57 S0:F127 s:F128 vdd:F129 vdds:F126 PSVTGP W=1.09u L=0.06u 
MMM57@2 S0:F133 s:F132 vdd:F131 vdds:F130 PSVTGP W=1.09u L=0.06u 
MMM58 CO:F135 co1:F136 vdd:F137 vdds:F134 PSVTGP W=1.09u L=0.06u 
MMM58@2 CO:F141 co1:F140 vdd:F139 vdds:F138 PSVTGP W=1.09u L=0.06u 
MMM59 CO:F75 co1:F76 gnd:F77 gnds:F74 NSVTGP W=0.77u L=0.06u 
MMM59@2 CO:F81 co1:F80 gnd:F79 gnds:F78 NSVTGP W=0.77u L=0.06u 
R1 axorb:F89 axorb:F116 171.028
R10 axorb:F60 axorb:F52 528.991
R100 s:F128 s:F121 656.025
R101 s:F128 s:F72 229.23
R102 s:F128 s:F68 81.0919
R103 s:F128 s:F61 658.597
R104 s:F132 s:F121 1854.45
R105 s:F132 s:F72 73.7117
R106 s:F132 s:F68 229.23
R107 s:F132 s:F61 1861.72
R108 s:F68 s:F121 388.756
R109 s:F68 s:F72 135.84
R11 axorb:F29 axorb:F23 0.001
R110 s:F68 s:F61 390.279
R111 s:F72 s:F121 1098.93
R112 s:F72 s:F61 1103.24
R113 s:F121 s:F115 0.001
R114 s:F121 s:F61 95.6383
R115 s:F61 s:F55 0.001
R116 CI CI:F5 0.001
R117 CI:F124 CI:F119 4149.35
R118 CI:F124 CI:F5 73.4079
R119 CI:F119 CI:F5 38.6696
R12 nb:F85 nb:F101 150.607
R120 CI:F5 CI:F64 60.5851
R121 CI:F5 CI:F59 39.7196
R122 CI:F59 CI:F64 2222.37
R123 gnd gnd:F8 0.001
R124 gnd:73 gnd:F8 6.20535
R125 gnd:73 gnd:371 8.17681
R126 gnd:F8 gnd:F79 40.8195
R127 gnd:F8 gnd:F77 40.6821
R128 gnd:F8 gnd:F69 40.8519
R129 gnd:F8 gnd:F39 38.8467
R13 nb:F85 nb:F41 157.906
R130 gnd:F8 gnd:371 7.70825
R131 gnd:F69 gnd:F79 1623.73
R132 gnd:F69 gnd:F77 1618.26
R133 gnd:F69 gnd:F63 0.001
R134 gnd:F69 gnd:F39 4386.57
R135 gnd:F77 gnd:F79 1616.98
R136 gnd:F77 gnd:F71 0.001
R137 gnd:F77 gnd:F39 4368.34
R138 gnd:F79 gnd:F39 4383.08
R139 gnd:F39 gnd:F45 0.001
R14 nb:F85 nb:F25 151.307
R140 vdd vdd:F10 0.001
R141 vdd:F10 vdd:F139 21.0201
R142 vdd:F10 vdd:F137 41.6097
R143 vdd:F10 vdd:F129 41.7843
R144 vdd:F10 vdd:F105 39.1857
R145 vdd:F129 vdd:F139 838.192
R146 vdd:F129 vdd:F137 1659.21
R147 vdd:F129 vdd:F123 0.001
R148 vdd:F129 vdd:F105 4408.16
R149 vdd:F137 vdd:F139 834.688
R15 nb:F101 nb:F95 0.001
R150 vdd:F137 vdd:F131 0.001
R151 vdd:F137 vdd:F105 4389.73
R152 vdd:F139 vdd:F105 2217.58
