
***Library file consisting only the library cell instances in the /pnr/op_data/b01_final_new.dspf file

***Library cell instances: 
***Total number of cell instances: 16
**HS65_GS_BFX284
**HS65_GS_DFPQX4
**HS65_GS_DFPQX9
**HS65_GS_NAND2X7
**HS65_GS_NOR4ABX2
**HS65_GS_NOR2X6
**HS65_GS_AOI22X6
**HS65_GS_AOI32X5
**HS65_GS_CBI4I6X5
**HS65_GS_OAI21X3
**HS65_GS_CB4I6X9
**HS65_GSS_XOR2X6
**HS65_GS_NOR2AX3
**HS65_GS_MUX21X4
**HS65_GS_AOI12X2
**HS65_GS_IVX9


.SUBCKT HS65_GSS_XOR2X6 Z B A gnd gnd vdd vdd
*modified
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 11:59 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.212 PJ=7.32
MMMN0 Z:F26 net60:F27 gnd gnd NSVTGP AD=0.0678255p AS=0.0820989p L=0.06u NRD=0.285714 NRS=0.261905 PD=0.254681u PS=0.742737u W=0.63u lpe=3 ngcon=1 po2act=0.295877 sca=3.79615 scb=0.00291824 scc=5.79832e-05
MMMN1 net60:F18 B:F19 gnd gnd NSVTGP AD=0.032p AS=0.0528p L=0.06u NRD=0.34375 NRS=0.34375 PD=0.2u PS=0.65u W=0.32u lpe=3 ngcon=1 po2act=0.260348 sca=12.7654 scb=0.014473 scc=0.00123392
MMMN2 net72:F36 A:F35 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.0585p as=0.1482p lpe=3 ngcon=1 nrd=0.0961538 nrs=0.358974 pd=0.15u po2act=0.288029 ps=1.16u sca=6.99142 scb=0.00671895 scc=0.000548722
MMMN3 Z:F32 B:F31 net72:F30 gnd NSVTGP L=0.06u W=0.78u ad=0.0839745p as=0.0585p lpe=3 ngcon=1 nrd=0.307692 nrs=0.0961538 pd=0.315319u po2act=0.357315 ps=0.15u sca=6.99117 scb=0.00671895 scc=0.000548722
MMMN4 net60:F24 A:F23 gnd gnd NSVTGP L=0.06u W=0.32u ad=0.032p as=0.0417011p lpe=3 ngcon=1 nrd=0.34375 nrs=0.407237 pd=0.2u po2act=0.311209 ps=0.377263u sca=12.765 scb=0.014473 scc=0.00123392
MMMP0 Z:F50 B:F51 net54:F52 vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=0.503896 sca=5.22195 scb=0.00477169 scc=0.000389094
MMMP1 net54:F46 net60:F47 vdd vdd PSVTGP AD=0.11p AS=0.1219p L=0.06u NRD=0.25 NRS=0.272727 PD=0.2u PS=0.693333u W=1.1u lpe=3 ngcon=1 po2act=0.358612 sca=5.22185 scb=0.00477169 scc=0.000389094
MMMP2 Z:F56 A:F55 net54:F54 vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.2145p lpe=3 ngcon=1 nrd=0.25 nrs=0.272727 pd=0.2u po2act=0.317336 ps=1.49u sca=5.22243 scb=0.00477169 scc=0.000389094
MMMP3 net60:F40 B:F39 net42:F38 vdd PSVTGP L=0.06u W=0.55u ad=0.099p as=0.045375p lpe=3 ngcon=1 nrd=0.3 nrs=0.15 pd=0.91u po2act=0.312353 ps=0.165u sca=5.35408 scb=0.00535557 scc=0.000199694
MMMP4 net42:F44 A:F43 vdd vdd PSVTGP L=0.06u W=0.55u ad=0.045375p as=0.06095p lpe=3 ngcon=1 nrd=0.15 nrs=0.201488 pd=0.165u po2act=0.568787 ps=0.346667u sca=5.35356 scb=0.00535557 scc=0.000199694
R1 gnd gnd 0.001
R10 Z:F50 Z:F5 38.5454
R11 Z:F5 Z:F26 38.2464
R12 Z:F26 Z:F32 0.001
R13 net54:F46 net54:F54 75.6297
R14 net54:F46 net54:F52 0.001
R15 B B:F4 0.001
R16 B:F51 B:F31 72.8046
R17 B:F51 B:F4 83.525
R18 B:F39 B:F19 110.552
R19 B:F39 B:F4 73.867
R2 gnd gnd 37.794
R20 B:F4 B:F31 133.242
R21 B:F4 B:F19 193.519
R22 net60:F47 net60:F40 256.621
R23 net60:F47 net60:F27 127.682
R24 net60:F47 net60:F18 248.978
R25 net60:F40 net60:F27 427.482
R26 net60:F40 net60:F18 100.946
R27 net60:F27 net60:F18 414.751
R28 net60:F18 net60:F24 0.001
R29 vdd vdd 0.001
R3 gnd gnd 37.9928
R30 vdd vdd 0.001
R31 vdd vdd 0.001
R32 vdd vdd 0.001
R33 vdd vdd 0.001
R34 vdd vdd 0.001
R35 vdd vdd 37.6272
R36 vdd vdd 0.001
R37 vdd vdd 37.623
R38 vdd vdd 0.001
R39 A A:F3 0.001
R4 gnd gnd 37.7205
R40 A:F3 A:F55 95.8674
R41 A:F3 A:F35 105.753
R42 A:F3 A:F23 61.2066
R43 A:F55 A:F35 68.2517
R44 A:F43 A:F23 98.7499
R45 gnd gnd 0.001
R46 gnd gnd 0.0256454
R47 gnd gnd 37.6237
R48 gnd gnd 0.001
R49 gnd gnd 0.001
R5 gnd gnd 0.001
R50 gnd gnd 0.001
R51 gnd gnd 0.001
R6 net42:F38 net42:F44 0.001
R7 net72:F30 net72:F36 0.001
R8 Z Z:F5 0.001
R9 Z:F50 Z:F56 0.001
.ENDS HS65_GSS_XOR2X6


.SUBCKT HS65_GS_AOI12X2 Z C B A gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:37 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=2.336 PJ=6.12
MMM43 Z:F31 B:F30 net036:F29 vdd PSVTGP L=0.06u W=0.31u ad=0.0867875p as=0.0562954p lpe=3 ngcon=1 nrd=4.63266 nrs=0.5858 pd=1.105u po2act=0.183784 ps=0.588041u sca=13.4931 scb=0.0152609 scc=0.00137372
MMM47 net036:F39 C:F38 vdd vdd PSVTGP L=0.06u W=0.35u ad=0.0635593p as=0.06125p lpe=3 ngcon=1 nrd=0.518851 nrs=0.314286 pd=0.663918u po2act=0.240634 ps=0.7u sca=1.21937 scb=3.09432e-05 scc=1.70794e-09
MMM52 Z:F35 A:F34 net036:F33 vdd PSVTGP L=0.06u W=0.31u ad=0.0867875p as=0.0562954p lpe=3 ngcon=1 nrd=2.32711 nrs=0.5858 pd=1.105u po2act=0.246559 ps=0.588041u sca=1.18857 scb=2.39069e-05 scc=9.01275e-10
MMM77 Z:F27 C:F26 gnd gnd NSVTGP L=0.06u W=0.205u ad=0.0216714p as=0.03485p lpe=3 ngcon=1 nrd=0.292683 nrs=0.268293 pd=0.205u po2act=0.268642 ps=0.545u sca=3.3841 scb=0.00192275 scc=8.55396e-06
MMM78 Z:F21 B:F22 net0134:F23 gnd NSVTGP AD=0.0264286p AS=0.018125p L=0.06u NRD=0.22 NRS=0.29 PD=0.25u PS=0.145u W=0.25u lpe=3 ngcon=1 po2act=0.339844 sca=3.20484 scb=0.00168506 scc=7.10806e-06
MMM79 net0134:F17 A:F18 gnd gnd NSVTGP AD=0.018125p AS=0.0425p L=0.06u NRD=0.29 NRS=0.22 PD=0.145u PS=0.59u W=0.25u lpe=3 ngcon=1 po2act=0.259976 sca=3.20494 scb=0.00168506 scc=7.10806e-06
R1 net0134:F17 net0134:F23 0.001
R10 net036:F33 net036:F29 0.001
R11 C C:F5 0.001
R12 C:F38 C:F26 1482.45
R13 C:F38 C:F5 200.161
R14 C:F5 C:F26 102.975
R15 A A:F3 0.001
R16 A:F34 A:F18 873.42
R17 A:F34 A:F3 1251.16
R18 A:F3 A:F18 66.4779
R19 Z Z:F6 0.001
R2 gnd gnd 0.001
R20 Z:F35 Z:F31 0.001
R21 Z:F35 Z:F6 38.9465
R22 Z:F6 Z:F21 38.3305
R23 Z:F21 Z:F27 0.001
R24 vdd vdd 0.001
R25 vdd vdd 0.001
R26 vdd vdd 0.001
R27 vdd vdd 0.001
R28 vdd vdd 37.6252
R29 vdd vdd 0.001
R3 gnd gnd 37.9283
R30 vdd vdd 37.685
R31 gnd gnd 0.001
R32 gnd gnd 0.0256454
R33 gnd gnd 37.6237
R34 gnd gnd 0.001
R35 gnd gnd 0.001
R4 gnd gnd 37.6765
R5 B B:F4 0.001
R6 B:F4 B:F30 73.5194
R7 B:F4 B:F22 285.562
R8 B:F30 B:F22 199.408
R9 net036:F33 net036:F39 0.001
.ENDS HS65_GS_AOI12X2


.SUBCKT HS65_GS_AOI12X23 Z C B A gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:37 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=5.84 PJ=10.92
MMM31 net0134:F47 A:F46 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.0804894p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=0.2u po2act=0.754548 ps=0.304255u sca=6.98478 scb=0.00671895 scc=0.000548722
MMM32 Z:F95 A:F94 net0116:F93 vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=1.50184 ps=0.2u sca=5.21258 scb=0.00477169 scc=0.000389094
MMM35 Z:F71 A:F70 net0116:F69 vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=0.739912 ps=0.2u sca=5.21474 scb=0.00477169 scc=0.000389094
MMM39 Z:F79 B:F78 net0116:F77 vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=1.33253 ps=0.2u sca=5.21304 scb=0.00477169 scc=0.000389094
MMM41 Z:F81 B:F82 net0116:F83 vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=1.50184 sca=5.21258 scb=0.00477169 scc=0.000389094
MMM42 Z:F87 B:F86 net0116:F85 vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=1.5865 ps=0.2u sca=5.21234 scb=0.00477169 scc=0.000389094
MMM43 Z:F89 B:F90 net0116:F91 vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=1.5865 sca=5.21234 scb=0.00477169 scc=0.000389094
MMM47 net0116:F101 C:F102 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=1.07856 sca=5.21376 scb=0.00477169 scc=0.000389094
MMM49 net0116:F107 C:F106 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=0.739912 ps=0.2u sca=5.21474 scb=0.00477169 scc=0.000389094
MMM52 Z:F65 A:F66 net0116:F67 vdd PSVTGP AD=0.11p AS=0.1838p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=1.45u W=1.1u lpe=3 ngcon=1 po2act=0.316529 sca=5.21602 scb=0.00477169 scc=0.000389094
MMM54 net0134:F23 A:F22 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=0.2u po2act=0.729259 ps=0.2u sca=6.9861 scb=0.00671895 scc=0.000548722
MMM57 net0134:F25 A:F26 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.282051 NRS=0.282051 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=1.04706 sca=6.98551 scb=0.00671895 scc=0.000548722
MMM58 Z:F29 B:F30 net0134:F31 gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.282051 NRS=0.282051 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=1.26703 sca=6.98507 scb=0.00671895 scc=0.000548722
MMM61 Z:F35 B:F34 net0134:F33 gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=0.2u po2act=1.38376 ps=0.2u sca=6.98478 scb=0.00671895 scc=0.000548722
MMM63 net0116:F109 C:F110 vdd vdd PSVTGP AD=0.1838p AS=0.11p L=0.06u NRD=0.25 NRS=0.25 PD=1.45u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=0.316529 sca=5.21602 scb=0.00477169 scc=0.000389094
MMM64 Z:F37 B:F38 net0134:F39 gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.282051 NRS=0.282051 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=1.38473 sca=6.98464 scb=0.00671895 scc=0.000548722
MMM65 net0116:F99 C:F98 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=1.33253 ps=0.2u sca=5.21304 scb=0.00477169 scc=0.000389094
MMM70 Z:F73 A:F74 net0116:F75 vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=1.07856 sca=5.21376 scb=0.00477169 scc=0.000389094
MMM73 Z:F63 C:F62 gnd gnd NSVTGP L=0.06u W=0.63u ad=0.063p as=0.10625p lpe=3 ngcon=1 nrd=0.261905 nrs=0.261905 pd=0.2u po2act=0.319267 ps=0.98u sca=3.79214 scb=0.00291824 scc=5.79832e-05
MMM75 Z:F49 C:F50 gnd gnd NSVTGP AD=0.063p AS=0.0650106p L=0.06u NRD=0.261905 NRS=0.261905 PD=0.2u PS=0.245745u W=0.63u lpe=3 ngcon=1 po2act=1.33434 sca=3.79014 scb=0.00291824 scc=5.79832e-05
MMM76 Z:F55 C:F54 gnd gnd NSVTGP L=0.06u W=0.63u ad=0.063p as=0.063p lpe=3 ngcon=1 nrd=0.261905 nrs=0.261905 pd=0.2u po2act=1.08061 ps=0.2u sca=3.79058 scb=0.00291824 scc=5.79832e-05
MMM77 Z:F57 C:F58 gnd gnd NSVTGP AD=0.063p AS=0.063p L=0.06u NRD=0.261905 NRS=0.261905 PD=0.2u PS=0.2u W=0.63u lpe=3 ngcon=1 po2act=0.742285 sca=3.79118 scb=0.00291824 scc=5.79832e-05
MMM78 Z:F43 B:F42 net0134:F41 gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=0.2u po2act=1.23321 ps=0.2u sca=6.98464 scb=0.00671895 scc=0.000548722
MMM79 net0134:F17 A:F18 gnd gnd NSVTGP AD=0.078p AS=0.131p L=0.06u NRD=0.282051 NRS=0.282051 PD=0.2u PS=1.13u W=0.78u lpe=3 ngcon=1 po2act=0.316266 sca=6.98706 scb=0.00671895 scc=0.000548722
R1 net0134:F17 net0134:F41 156.499
R10 net0134:F41 net0134:F47 0.001
R100 B:F90 B:F42 83.9431
R101 B:F90 B:F38 355.389
R102 B:F90 B:F34 1491.08
R103 B:F90 B:F30 4037.97
R104 B:F90 B:F4 188.135
R105 B:F4 B:F42 206.052
R106 B:F4 B:F38 190.537
R107 B:F4 B:F34 146.677
R108 B:F4 B:F30 397.212
R109 B:F38 B:F42 389.235
R11 Z Z:F6 0.001
R110 B:F38 B:F34 482.781
R111 B:F38 B:F30 1307.41
R112 B:F42 B:F34 1633.09
R113 B:F42 B:F30 4422.53
R114 B:F30 B:F34 347.744
R115 A A:F3 0.001
R116 A:F66 A:F74 1149.79
R117 A:F66 A:F70 332.417
R118 A:F66 A:F26 1259.29
R119 A:F66 A:F22 364.076
R12 Z:F57 Z:F63 0.001
R120 A:F66 A:F18 87.3444
R121 A:F66 A:F3 149.516
R122 A:F70 A:F74 332.358
R123 A:F70 A:F26 364.011
R124 A:F70 A:F22 105.24
R125 A:F70 A:F18 364.076
R126 A:F70 A:F3 149.809
R127 A:F22 A:F74 364.011
R128 A:F22 A:F26 398.679
R129 A:F22 A:F18 398.75
R13 Z:F57 Z:F49 2544.76
R130 A:F22 A:F3 164.076
R131 A:F74 A:F26 86.9923
R132 A:F74 A:F18 1259.29
R133 A:F74 A:F3 151.742
R134 A:F94 A:F46 69.6056
R135 A:F94 A:F3 111.902
R136 A:F3 A:F46 101.729
R137 A:F3 A:F26 166.194
R138 A:F3 A:F18 163.755
R139 A:F18 A:F26 1379.22
R14 Z:F57 Z:F37 2674.28
R140 vdd vdd 0.001
R141 vdd vdd 38.7875
R142 vdd vdd 38.657
R143 vdd vdd 0.001
R144 vdd vdd 2510.21
R145 vdd vdd 0.001
R146 vdd vdd 0.001
R147 vdd vdd 0.001
R148 vdd vdd 0.001
R149 vdd vdd 0.001
R15 Z:F57 Z:F29 2723.03
R150 vdd vdd 0.001
R151 vdd vdd 0.001
R152 vdd vdd 0.001
R153 vdd vdd 0.001
R154 vdd vdd 0.001
R155 vdd vdd 0.001
R156 vdd vdd 0.001
R157 vdd vdd 0.001
R158 vdd vdd 0.001
R159 vdd vdd 37.6252
R16 Z:F57 Z:F6 40.4834
R160 gnd gnd 0.001
R161 gnd gnd 0.0256454
R162 gnd gnd 37.6237
R163 gnd gnd 0.001
R164 gnd gnd 0.001
R165 gnd gnd 0.001
R166 gnd gnd 0.001
R167 gnd gnd 0.001
R168 gnd gnd 0.001
R169 gnd gnd 0.001
R17 Z:F71 Z:F95 2721.55
R170 gnd gnd 0.001
R171 gnd gnd 0.001
R172 gnd gnd 0.001
R173 gnd gnd 0.001
R174 C C:F5 0.001
R175 C:F5 C:F110 84.9896
R176 C:F5 C:F106 99.904
R177 C:F5 C:F102 271.528
R178 C:F5 C:F98 623.563
R179 C:F5 C:F62 214.497
R18 Z:F71 Z:F87 1351.53
R180 C:F5 C:F58 252.139
R181 C:F5 C:F54 685.285
R182 C:F5 C:F50 1573.76
R183 C:F50 C:F110 4279.54
R184 C:F50 C:F106 1464.75
R185 C:F50 C:F102 430.284
R186 C:F50 C:F98 140.542
R187 C:F50 C:F62 10800.7
R188 C:F50 C:F58 3696.75
R189 C:F50 C:F54 1085.95
R19 Z:F71 Z:F79 883.251
R190 C:F54 C:F110 1863.51
R191 C:F54 C:F106 637.82
R192 C:F54 C:F102 187.365
R193 C:F54 C:F98 430.284
R194 C:F54 C:F62 4703.14
R195 C:F54 C:F58 1609.74
R196 C:F58 C:F110 685.645
R197 C:F58 C:F106 234.675
R198 C:F58 C:F102 637.82
R199 C:F58 C:F98 1464.75
R2 net0134:F17 net0134:F33 153.86
R20 Z:F71 Z:F65 0.001
R200 C:F58 C:F62 1730.44
R201 C:F98 C:F110 1695.67
R202 C:F98 C:F106 580.373
R203 C:F98 C:F102 170.49
R204 C:F98 C:F62 4279.54
R205 C:F102 C:F110 738.371
R206 C:F102 C:F106 252.721
R207 C:F102 C:F62 1863.51
R208 C:F106 C:F110 271.67
R209 C:F106 C:F62 685.644
R21 Z:F71 Z:F6 43.6669
R210 C:F110 C:F62 190.731
R22 Z:F79 Z:F95 2664.75
R23 Z:F79 Z:F87 1622.41
R24 Z:F79 Z:F73 0.001
R25 Z:F79 Z:F6 42.7556
R26 Z:F87 Z:F95 2595.79
R27 Z:F87 Z:F81 0.001
R28 Z:F87 Z:F6 41.6491
R29 Z:F95 Z:F89 0.001
R3 net0134:F17 net0134:F25 148.798
R30 Z:F95 Z:F6 39.7845
R31 Z:F6 Z:F49 39.8084
R32 Z:F6 Z:F37 41.8345
R33 Z:F6 Z:F29 42.597
R34 Z:F29 Z:F49 2677.62
R35 Z:F29 Z:F37 1004.73
R36 Z:F29 Z:F35 0.001
R37 Z:F37 Z:F49 2629.69
R38 Z:F37 Z:F43 0.001
R39 Z:F49 Z:F55 0.001
R4 net0134:F17 net0134:F23 0.001
R40 gnd gnd 0.001
R41 gnd gnd 2359.52
R42 gnd gnd 0.001
R43 gnd gnd 2357.92
R44 gnd gnd 39.3802
R45 gnd gnd 39.5131
R46 gnd gnd 39.4862
R47 gnd gnd 37.5904
R48 gnd gnd 37.5
R49 gnd gnd 2365.88
R5 net0134:F25 net0134:F41 153.86
R50 gnd gnd 0.001
R51 gnd gnd 0.001
R52 net0116:F107 net0116:F109 239.634
R53 net0116:F107 net0116:F101 0.001
R54 net0116:F107 net0116:F99 252.2
R55 net0116:F107 net0116:F91 266.375
R56 net0116:F107 net0116:F83 277.892
R57 net0116:F107 net0116:F75 286.036
R58 net0116:F107 net0116:F67 290.258
R59 net0116:F109 net0116:F99 255.923
R6 net0134:F25 net0134:F33 151.265
R60 net0116:F109 net0116:F91 270.307
R61 net0116:F109 net0116:F83 281.994
R62 net0116:F109 net0116:F75 290.258
R63 net0116:F109 net0116:F67 294.543
R64 net0116:F99 net0116:F93 0.001
R65 net0116:F99 net0116:F91 258.79
R66 net0116:F99 net0116:F83 269.979
R67 net0116:F99 net0116:F75 277.892
R68 net0116:F99 net0116:F67 281.994
R69 net0116:F67 net0116:F91 270.307
R7 net0134:F25 net0134:F31 0.001
R70 net0116:F67 net0116:F83 255.923
R71 net0116:F67 net0116:F75 239.634
R72 net0116:F75 net0116:F91 266.375
R73 net0116:F75 net0116:F83 252.2
R74 net0116:F75 net0116:F69 0.001
R75 net0116:F83 net0116:F91 258.79
R76 net0116:F83 net0116:F77 0.001
R77 net0116:F91 net0116:F85 0.001
R78 B B:F4 0.001
R79 B:F86 B:F90 324.485
R8 net0134:F33 net0134:F41 148.798
R80 B:F86 B:F82 402.47
R81 B:F86 B:F78 1089.92
R82 B:F86 B:F42 355.389
R83 B:F86 B:F38 105.061
R84 B:F86 B:F34 440.8
R85 B:F86 B:F30 1193.72
R86 B:F86 B:F4 173.968
R87 B:F78 B:F90 3686.84
R88 B:F78 B:F82 289.896
R89 B:F78 B:F42 4037.97
R9 net0134:F33 net0134:F39 0.001
R90 B:F78 B:F38 1193.72
R91 B:F78 B:F34 317.505
R92 B:F78 B:F30 79.1708
R93 B:F78 B:F4 362.672
R94 B:F82 B:F90 1361.42
R95 B:F82 B:F42 1491.08
R96 B:F82 B:F38 440.8
R97 B:F82 B:F34 117.244
R98 B:F82 B:F30 317.506
R99 B:F82 B:F4 133.922
.ENDS HS65_GS_AOI12X23


.SUBCKT HS65_GS_AOI22X6 Z D C B A gnd gnd vdd vdd
*MOdified
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:08 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=2.92 PJ=6.92
MMM12 net0161:F33 A:F32 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.0663p as=0.1755p lpe=3 ngcon=1 nrd=0.108974 nrs=0.410256 pd=0.17u po2act=0.365625 ps=1.23u sca=6.99217 scb=0.00671895 scc=0.000548722
MMM13 net0244:F47 A:F48 vdd vdd PSVTGP AD=0.22p AS=0.121p L=0.06u NRD=0.272727 NRS=0.295455 PD=1.5u PS=0.22u W=1.1u lpe=3 ngcon=1 po2act=0.333884 sca=5.22363 scb=0.00477169 scc=0.000389094
MMM15 net0244:F45 B:F44 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.1155p as=0.121p lpe=3 ngcon=1 nrd=0.272727 nrs=0.295455 pd=0.21u po2act=0.579174 ps=0.22u sca=5.22318 scb=0.00477169 scc=0.000389094
MMM16 Z:F35 C:F36 net0244:F37 vdd PSVTGP AD=0.1155p AS=0.209p L=0.06u NRD=0.272727 NRS=0.272727 PD=0.21u PS=1.48u W=1.1u lpe=3 ngcon=1 po2act=0.320331 sca=5.22365 scb=0.00477169 scc=0.000389094
MMM17 Z:F41 D:F40 net0244:F39 vdd PSVTGP L=0.06u W=1.1u ad=0.1155p as=0.1155p lpe=3 ngcon=1 nrd=0.272727 nrs=0.272727 pd=0.21u po2act=0.570248 ps=0.21u sca=5.2232 scb=0.00477169 scc=0.000389094
MMM23 Z:F23 D:F24 net038:F25 gnd NSVTGP AD=0.0858p AS=0.08385p L=0.06u NRD=0.333333 NRS=0.137821 PD=0.22u PS=0.215u W=0.78u lpe=3 ngcon=1 po2act=0.569625 sca=6.99197 scb=0.00671895 scc=0.000548722
MMM24 net038:F19 C:F20 gnd gnd NSVTGP AD=0.08385p AS=0.1482p L=0.06u NRD=0.137821 NRS=0.307692 PD=0.215u PS=1.16u W=0.78u lpe=3 ngcon=1 po2act=0.319833 sca=6.99223 scb=0.00671895 scc=0.000548722
MMM8 Z:F29 B:F28 net0161:F27 gnd NSVTGP L=0.06u W=0.78u ad=0.0858p as=0.0663p lpe=3 ngcon=1 nrd=0.333333 nrs=0.108974 pd=0.22u po2act=0.564958 ps=0.17u sca=6.99197 scb=0.00671895 scc=0.000548722
R1 net0161:F27 net0161:F33 0.001
R10 Z Z:F7 0.001
R11 Z:F41 Z:F35 0.001
R12 Z:F41 Z:F7 37.6912
R13 Z:F7 Z:F23 39.7243
R14 Z:F23 Z:F29 0.001
R15 B B:F4 0.001
R16 B:F44 B:F28 72.3727
R17 B:F44 B:F4 102.122
R18 B:F4 B:F28 102.122
R19 D D:F6 0.001
R2 net038:F19 net038:F25 0.001
R20 D:F40 D:F24 74.264
R21 D:F40 D:F6 102.393
R22 D:F6 D:F24 102.393
R23 C C:F5 0.001
R24 C:F36 C:F5 100.244
R25 C:F36 C:F20 66.5044
R26 C:F5 C:F20 100.244
R27 net0244:F37 net0244:F47 114.83
R28 net0244:F37 net0244:F39 113.064
R29 net0244:F39 net0244:F47 113.096
R3 gnd gnd 0.001
R30 net0244:F39 net0244:F45 0.001
R31 vdd vdd 0.001
R32 vdd vdd 0.001
R33 vdd vdd 0.001
R34 vdd vdd 0.001
R35 vdd vdd 0.001
R36 vdd vdd 37.6252
R37 vdd vdd 0.001
R38 vdd vdd 37.7106
R39 vdd vdd 0.001
R4 gnd gnd 37.5373
R40 gnd gnd 0.001
R41 gnd gnd 0.001
R42 gnd gnd 0.001
R43 gnd gnd 0.001
R44 gnd gnd 0.0256454
R45 gnd gnd 37.6237
R5 gnd gnd 37.7737
R6 A A:F3 0.001
R7 A:F48 A:F32 67.4722
R8 A:F48 A:F3 118.295
R9 A:F3 A:F32 118.295
.ENDS HS65_GS_AOI22X6


.SUBCKT HS65_GS_AOI32X5 Z E D C B A gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:09 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.212 PJ=7.32
MMM10 net0161:F35 B:F34 net034:F33 gnd NSVTGP L=0.06u W=0.78u ad=0.07215p as=0.07215p lpe=3 ngcon=1 nrd=0.11859 nrs=0.11859 pd=0.185u po2act=0.623298 ps=0.185u sca=6.99117 scb=0.00671895 scc=0.000548722
MMM12 net034:F39 A:F38 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.07215p as=0.1716p lpe=3 ngcon=1 nrd=0.11859 nrs=0.410256 pd=0.185u po2act=0.371348 ps=1.22u sca=6.99146 scb=0.00671895 scc=0.000548722
MMM13 net0244:F59 A:F58 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.1155p as=0.198p lpe=3 ngcon=1 nrd=0.272727 nrs=0.272727 pd=0.21u po2act=0.314043 ps=1.46u sca=5.22262 scb=0.00477169 scc=0.000389094
MMM15 net0244:F51 C:F50 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=0.704965 ps=0.2u sca=5.22184 scb=0.00477169 scc=0.000389094
MMM16 Z:F41 D:F42 net0244:F43 vdd PSVTGP AD=0.11p AS=0.198p L=0.06u NRD=0.25 NRS=0.272727 PD=0.2u PS=1.46u W=1.1u lpe=3 ngcon=1 po2act=0.314043 sca=5.22262 scb=0.00477169 scc=0.000389094
MMM22 net029:F21 D:F22 gnd gnd NSVTGP AD=0.06435p AS=0.1404p L=0.06u NRD=0.105769 NRS=0.307692 PD=0.165u PS=1.14u W=0.78u lpe=3 ngcon=1 po2act=0.314043 sca=6.99152 scb=0.00671895 scc=0.000548722
MMM23 Z:F25 E:F26 net029:F27 gnd NSVTGP AD=0.09165p AS=0.06435p L=0.06u NRD=0.384615 NRS=0.105769 PD=0.235u PS=0.165u W=0.78u lpe=3 ngcon=1 po2act=0.57734 sca=6.99122 scb=0.00671895 scc=0.000548722
MMM27 Z:F47 E:F46 net0244:F45 vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=0.60539 ps=0.2u sca=5.22203 scb=0.00477169 scc=0.000389094
MMM28 net0244:F53 B:F54 vdd vdd PSVTGP AD=0.1155p AS=0.11p L=0.06u NRD=0.272727 NRS=0.25 PD=0.21u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=0.612766 sca=5.22202 scb=0.00477169 scc=0.000389094
MMM8 Z:F31 C:F30 net0161:F29 gnd NSVTGP L=0.06u W=0.78u ad=0.09165p as=0.07215p lpe=3 ngcon=1 nrd=0.358974 nrs=0.11859 pd=0.235u po2act=0.704965 ps=0.185u sca=6.99107 scb=0.00671895 scc=0.000548722
R1 net034:F33 net034:F39 0.001
R10 A:F3 A:F38 99.0743
R11 B B:F4 0.001
R12 B:F54 B:F4 103.037
R13 B:F54 B:F34 76.3586
R14 B:F4 B:F34 103.037
R15 Z Z:F8 0.001
R16 Z:F47 Z:F41 0.001
R17 Z:F47 Z:F8 38.2626
R18 Z:F8 Z:F25 39.7965
R19 Z:F25 Z:F31 0.001
R2 net0161:F29 net0161:F35 0.001
R20 C C:F5 0.001
R21 C:F50 C:F5 103.711
R22 C:F50 C:F30 77.4419
R23 C:F5 C:F30 103.711
R24 E E:F7 0.001
R25 E:F46 E:F7 103.243
R26 E:F46 E:F26 76.3023
R27 E:F7 E:F26 103.243
R28 D D:F6 0.001
R29 D:F42 D:F6 101.771
R3 net029:F21 net029:F27 0.001
R30 D:F42 D:F22 70.7482
R31 D:F6 D:F22 101.771
R32 net0244:F43 net0244:F53 115.233
R33 net0244:F43 net0244:F45 113.18
R34 net0244:F45 net0244:F53 113.18
R35 net0244:F45 net0244:F51 0.001
R36 net0244:F53 net0244:F59 0.001
R37 vdd vdd 0.001
R38 vdd vdd 0.001
R39 vdd vdd 0.001
R4 gnd gnd 0.001
R40 vdd vdd 0.001
R41 vdd vdd 0.001
R42 vdd vdd 0.001
R43 vdd vdd 37.6252
R44 vdd vdd 0.001
R45 vdd vdd 37.8301
R46 vdd vdd 37.901
R47 vdd vdd 0.001
R48 gnd gnd 0.001
R49 gnd gnd 0.001
R5 gnd gnd 37.5
R50 gnd gnd 0.001
R51 gnd gnd 0.001
R52 gnd gnd 0.001
R53 gnd gnd 0.0256454
R54 gnd gnd 37.6237
R6 gnd gnd 37.8086
R7 A A:F3 0.001
R8 A:F58 A:F38 63.1849
R9 A:F58 A:F3 99.0743
.ENDS HS65_GS_AOI32X5


.SUBCKT HS65_GS_BFX284 Z A gnd gnd vdd vdd

*Modified subckt

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:10 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=17.812 PJ=27.32
MMM0 net0513:F142 A:F143 gnd gnd NSVTGP AD=0.0819p AS=0.078p L=0.06u NRD=0.153846 NRS=0.141026 PD=0.21u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=4.34057 sca=6.97812 scb=0.00671895 scc=0.000548722
MMM1 net0513:F148 A:F147 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.0819p as=0.0819p lpe=3 ngcon=1 nrd=0.153846 nrs=0.153846 pd=0.21u po2act=4.0637 ps=0.21u sca=6.97868 scb=0.00671895 scc=0.000548722
MMM10 net0513:F182 A:F183 gnd gnd NSVTGP AD=0.1521p AS=0.0897p L=0.06u NRD=0.179487 NRS=0.179487 PD=1.17u PS=0.23u W=0.78u lpe=3 ngcon=1 po2act=0.38254 sca=6.98696 scb=0.00671895 scc=0.000548722
MMM11 net0513:F314 A:F315 vdd vdd PSVTGP AD=0.1155p AS=0.11p L=0.06u NRD=0.136364 NRS=0.125 PD=0.21u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=4.34057 sca=5.20084 scb=0.00477169 scc=0.000389094
MMM12 net0513:F320 A:F319 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.1155p as=0.1155p lpe=3 ngcon=1 nrd=0.136364 nrs=0.136364 pd=0.21u po2act=4.0637 ps=0.21u sca=5.20161 scb=0.00477169 scc=0.000389094
MMM13 net0513:F322 A:F323 vdd vdd PSVTGP AD=0.1155p AS=0.1155p L=0.06u NRD=0.136364 NRS=0.136364 PD=0.21u PS=0.21u W=1.1u lpe=3 ngcon=1 po2act=3.76128 sca=5.20246 scb=0.00477169 scc=0.000389094
MMM14 net0513:F328 A:F327 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.1155p as=0.1155p lpe=3 ngcon=1 nrd=0.136364 nrs=0.136364 pd=0.21u po2act=3.43331 ps=0.21u sca=5.20339 scb=0.00477169 scc=0.000389094
MMM15 net0513:F330 A:F331 vdd vdd PSVTGP AD=0.1155p AS=0.1155p L=0.06u NRD=0.136364 NRS=0.136364 PD=0.21u PS=0.21u W=1.1u lpe=3 ngcon=1 po2act=3.07978 sca=5.20442 scb=0.00477169 scc=0.000389094
MMM16 net0513:F336 A:F335 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.1155p as=0.1155p lpe=3 ngcon=1 nrd=0.136364 nrs=0.136364 pd=0.21u po2act=2.70069 ps=0.21u sca=5.20557 scb=0.00477169 scc=0.000389094
MMM17 net0513:F338 A:F339 vdd vdd PSVTGP AD=0.1155p AS=0.1155p L=0.06u NRD=0.136364 NRS=0.136364 PD=0.21u PS=0.21u W=1.1u lpe=3 ngcon=1 po2act=2.29305 sca=5.20683 scb=0.00477169 scc=0.000389094
MMM18 net0513:F344 A:F343 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.1155p as=0.1155p lpe=3 ngcon=1 nrd=0.136364 nrs=0.136364 pd=0.21u po2act=1.85941 ps=0.21u sca=5.20825 scb=0.00477169 scc=0.000389094
MMM19 net0513:F346 A:F347 vdd vdd PSVTGP AD=0.1155p AS=0.1155p L=0.06u NRD=0.136364 NRS=0.136364 PD=0.21u PS=0.21u W=1.1u lpe=3 ngcon=1 po2act=1.404 sca=5.20983 scb=0.00477169 scc=0.000389094
MMM2 net0513:F150 A:F151 gnd gnd NSVTGP AD=0.0819p AS=0.0819p L=0.06u NRD=0.153846 NRS=0.153846 PD=0.21u PS=0.21u W=0.78u lpe=3 ngcon=1 po2act=3.76128 sca=6.97929 scb=0.00671895 scc=0.000548722
MMM20 net0513:F352 A:F351 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.1155p as=0.1265p lpe=3 ngcon=1 nrd=0.136364 nrs=0.159091 pd=0.21u po2act=0.925131 ps=0.23u sca=5.21162 scb=0.00477169 scc=0.000389094
MMM21 net0513:F354 A:F355 vdd vdd PSVTGP AD=0.2145p AS=0.1265p L=0.06u NRD=0.159091 NRS=0.159091 PD=1.49u PS=0.23u W=1.1u lpe=3 ngcon=1 po2act=0.38254 sca=5.2138 scb=0.00477169 scc=0.000389094
MMM3 net0513:F156 A:F155 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.0819p as=0.0819p lpe=3 ngcon=1 nrd=0.153846 nrs=0.153846 pd=0.21u po2act=3.43331 ps=0.21u sca=6.97995 scb=0.00671895 scc=0.000548722
MMM4 net0513:F158 A:F159 gnd gnd NSVTGP AD=0.0819p AS=0.0819p L=0.06u NRD=0.153846 NRS=0.153846 PD=0.21u PS=0.21u W=0.78u lpe=3 ngcon=1 po2act=3.07978 sca=6.98068 scb=0.00671895 scc=0.000548722
MMM5 net0513:F164 A:F163 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.0819p as=0.0819p lpe=3 ngcon=1 nrd=0.153846 nrs=0.153846 pd=0.21u po2act=2.70069 ps=0.21u sca=6.98147 scb=0.00671895 scc=0.000548722
MMM6 net0513:F166 A:F167 gnd gnd NSVTGP AD=0.0819p AS=0.0819p L=0.06u NRD=0.153846 NRS=0.153846 PD=0.21u PS=0.21u W=0.78u lpe=3 ngcon=1 po2act=2.29305 sca=6.98235 scb=0.00671895 scc=0.000548722
MMM7 net0513:F172 A:F171 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.0819p as=0.0819p lpe=3 ngcon=1 nrd=0.153846 nrs=0.153846 pd=0.21u po2act=1.85941 ps=0.21u sca=6.98331 scb=0.00671895 scc=0.000548722
MMM8 net0513:F174 A:F175 gnd gnd NSVTGP AD=0.0819p AS=0.0819p L=0.06u NRD=0.153846 NRS=0.153846 PD=0.21u PS=0.21u W=0.78u lpe=3 ngcon=1 po2act=1.404 sca=6.98437 scb=0.00671895 scc=0.000548722
MMM9 net0513:F180 A:F179 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.0819p as=0.0897p lpe=3 ngcon=1 nrd=0.153846 nrs=0.179487 pd=0.21u po2act=0.925131 ps=0.23u sca=6.98554 scb=0.00671895 scc=0.000548722
MMMI0 Z:F140 net0513:F139 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=4.58302 ps=0.2u sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI1 Z:F134 net0513:F135 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=4.80177 sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI10 Z:F100 net0513:F99 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=5.70414 ps=0.2u sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI11 Z:F94 net0513:F95 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=5.68591 sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI12 Z:F92 net0513:F91 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=5.64398 ps=0.2u sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI13 Z:F86 net0513:F87 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=5.57836 sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI14 Z:F84 net0513:F83 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=5.48903 ps=0.2u sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI15 Z:F78 net0513:F79 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=5.37601 sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI16 Z:F76 net0513:F75 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=5.23929 ps=0.2u sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI17 Z:F70 net0513:F71 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=5.07887 sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI18 Z:F68 net0513:F67 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=4.89475 ps=0.2u sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI19 Z:F62 net0513:F63 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=4.68693 sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI2 Z:F132 net0513:F131 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=4.99683 ps=0.2u sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI20 Z:F60 net0513:F59 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=4.45541 ps=0.2u sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI21 Z:F54 net0513:F55 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=4.2002 sca=6.9784 scb=0.00671895 scc=0.000548722
MMMI22 Z:F52 net0513:F51 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=3.92128 ps=0.2u sca=6.97897 scb=0.00671895 scc=0.000548722
MMMI23 Z:F46 net0513:F47 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=3.61867 sca=6.97958 scb=0.00671895 scc=0.000548722
MMMI24 Z:F44 net0513:F43 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=3.29236 ps=0.2u sca=6.98024 scb=0.00671895 scc=0.000548722
MMMI25 Z:F38 net0513:F39 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=2.94235 sca=6.98096 scb=0.00671895 scc=0.000548722
MMMI26 Z:F36 net0513:F35 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=2.56865 ps=0.2u sca=6.98175 scb=0.00671895 scc=0.000548722
MMMI27 Z:F30 net0513:F31 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=2.16674 sca=6.98262 scb=0.00671895 scc=0.000548722
MMMI28 Z:F28 net0513:F27 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=1.7435 ps=0.2u sca=6.98357 scb=0.00671895 scc=0.000548722
MMMI29 Z:F22 net0513:F23 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=1.29967 sca=6.98462 scb=0.00671895 scc=0.000548722
MMMI3 Z:F126 net0513:F127 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=5.16819 sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI30 Z:F20 net0513:F19 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=0.833733 ps=0.2u sca=6.98578 scb=0.00671895 scc=0.000548722
MMMI31 Z:F14 net0513:F15 gnd gnd NSVTGP AD=0.078p AS=0.1365p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=1.13u W=0.78u lpe=3 ngcon=1 po2act=0.34398 sca=6.98706 scb=0.00671895 scc=0.000548722
MMMI32 Z:F312 net0513:F311 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=4.58302 ps=0.2u sca=5.20016 scb=0.00477169 scc=0.000389094
MMMI33 Z:F306 net0513:F307 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=4.80177 sca=5.19953 scb=0.00477169 scc=0.000389094
MMMI34 Z:F304 net0513:F303 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=4.99683 ps=0.2u sca=5.19896 scb=0.00477169 scc=0.000389094
MMMI35 Z:F298 net0513:F299 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=5.16819 sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI36 Z:F296 net0513:F295 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=5.31585 ps=0.2u sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI37 Z:F290 net0513:F291 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=5.43981 sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI38 Z:F288 net0513:F287 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=5.54007 ps=0.2u sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI39 Z:F282 net0513:F283 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=5.61664 sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI4 Z:F124 net0513:F123 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=5.31585 ps=0.2u sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI40 Z:F280 net0513:F279 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=5.6695 ps=0.2u sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI41 Z:F274 net0513:F275 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=5.69867 sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI42 Z:F272 net0513:F271 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=5.70414 ps=0.2u sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI43 Z:F266 net0513:F267 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=5.68591 sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI44 Z:F264 net0513:F263 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=5.64398 ps=0.2u sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI45 Z:F258 net0513:F259 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=5.57836 sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI46 Z:F256 net0513:F255 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=5.48903 ps=0.2u sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI47 Z:F250 net0513:F251 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=5.37601 sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI48 Z:F248 net0513:F247 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=5.23929 ps=0.2u sca=5.19846 scb=0.00477169 scc=0.000389094
MMMI49 Z:F242 net0513:F243 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=5.07887 sca=5.1987 scb=0.00477169 scc=0.000389094
MMMI5 Z:F118 net0513:F119 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=5.43981 sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI50 Z:F240 net0513:F239 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=4.89475 ps=0.2u sca=5.19926 scb=0.00477169 scc=0.000389094
MMMI51 Z:F234 net0513:F235 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=4.68693 sca=5.19986 scb=0.00477169 scc=0.000389094
MMMI52 Z:F232 net0513:F231 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=4.45541 ps=0.2u sca=5.20052 scb=0.00477169 scc=0.000389094
MMMI53 Z:F226 net0513:F227 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=4.2002 sca=5.20123 scb=0.00477169 scc=0.000389094
MMMI54 Z:F224 net0513:F223 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=3.92128 ps=0.2u sca=5.20201 scb=0.00477169 scc=0.000389094
MMMI55 Z:F218 net0513:F219 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=3.61867 sca=5.20286 scb=0.00477169 scc=0.000389094
MMMI56 Z:F216 net0513:F215 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=3.29236 ps=0.2u sca=5.2038 scb=0.00477169 scc=0.000389094
MMMI57 Z:F210 net0513:F211 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=2.94235 sca=5.20483 scb=0.00477169 scc=0.000389094
MMMI58 Z:F208 net0513:F207 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=2.56865 ps=0.2u sca=5.20597 scb=0.00477169 scc=0.000389094
MMMI59 Z:F202 net0513:F203 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=2.16674 sca=5.20724 scb=0.00477169 scc=0.000389094
MMMI6 Z:F116 net0513:F115 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=5.54007 ps=0.2u sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI60 Z:F200 net0513:F199 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=1.7435 ps=0.2u sca=5.20864 scb=0.00477169 scc=0.000389094
MMMI61 Z:F194 net0513:F195 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=1.29967 sca=5.21021 scb=0.00477169 scc=0.000389094
MMMI62 Z:F192 net0513:F191 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.125 pd=0.2u po2act=0.833733 ps=0.2u sca=5.21197 scb=0.00477169 scc=0.000389094
MMMI63 Z:F186 net0513:F187 vdd vdd PSVTGP AD=0.11p AS=0.1925p L=0.06u NRD=0.125 NRS=0.125 PD=0.2u PS=1.45u W=1.1u lpe=3 ngcon=1 po2act=0.34398 sca=5.21396 scb=0.00477169 scc=0.000389094
MMMI7 Z:F110 net0513:F111 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=5.61664 sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI8 Z:F108 net0513:F107 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.141026 pd=0.2u po2act=5.6695 ps=0.2u sca=6.97808 scb=0.00671895 scc=0.000548722
MMMI9 Z:F102 net0513:F103 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.141026 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=5.69867 sca=6.97808 scb=0.00671895 scc=0.000548722
R1 vdd vdd 0.001
R10 vdd vdd 0.001
R100 A:F167 A:F171 513.088
R1000 net0513:F203 net0513:F15 11904
R1001 vdd vdd 0.001
R1002 vdd vdd 19.6053
R1003 vdd vdd 19.4667
R1004 vdd vdd 19.1536
R1005 vdd vdd 18.8094
R1006 vdd vdd 21.6499
R1007 vdd vdd 25.2053
R1008 vdd vdd 29.8872
R1009 vdd vdd 36.3039
R101 A:F167 A:F155 6679.64
R1010 vdd vdd 45.7604
R1011 vdd vdd 61.5944
R1012 vdd vdd 92.9095
R1013 vdd vdd 186.444
R1014 vdd vdd 1.25491
R1015 vdd vdd 179.539
R1016 vdd vdd 89.5725
R1017 vdd vdd 60.2317
R1018 vdd vdd 43.0553
R1019 vdd vdd 35.2701
R102 A:F167 A:F3 202.091
R1020 vdd vdd 29.5395
R1021 vdd vdd 24.6385
R1022 vdd vdd 21.083
R1023 vdd vdd 18.8094
R1024 vdd vdd 21.5552
R1025 vdd vdd 24.9953
R1026 vdd vdd 29.6374
R1027 vdd vdd 36.0004
R1028 vdd vdd 45.3779
R1029 vdd vdd 61.0795
R103 A:F171 A:F355 5599.46
R1030 vdd vdd 92.1328
R1031 vdd vdd 184.886
R1032 vdd vdd 1.24442
R1033 vdd vdd 160.452
R1034 vdd vdd 91.8248
R1035 vdd vdd 61.0795
R1036 vdd vdd 43.4249
R1037 vdd vdd 35.4583
R1038 vdd vdd 29.6374
R1039 vdd vdd 24.6836
R104 A:F171 A:F351 1604.81
R1040 vdd vdd 21.1031
R1041 vdd vdd 18.8134
R1042 vdd vdd 1176.64
R1043 vdd vdd 1170.04
R1044 vdd vdd 0.001
R1045 vdd vdd 880.061
R1046 vdd vdd 938.875
R1047 vdd vdd 1123.4
R1048 vdd vdd 0.001
R1049 vdd vdd 0.001
R105 A:F171 A:F347 490.301
R1050 vdd vdd 0.001
R1051 vdd vdd 1691.04
R1052 vdd vdd 0.001
R1053 vdd vdd 1397.58
R1054 vdd vdd 0.001
R1055 vdd vdd 0.001
R1056 vdd vdd 0.001
R1057 vdd vdd 0.001
R1058 vdd vdd 0.001
R1059 vdd vdd 1199.46
R106 A:F171 A:F343 105.689
R1060 vdd vdd 0.001
R1061 vdd vdd 895.053
R1062 vdd vdd 954.291
R1063 vdd vdd 1142.78
R1064 vdd vdd 0.001
R1065 vdd vdd 0.001
R1066 vdd vdd 0.001
R1067 vdd vdd 0.001
R1068 vdd vdd 0.001
R1069 vdd vdd 0.001
R107 A:F171 A:F339 446.164
R1070 vdd vdd 0.001
R1071 vdd vdd 0.001
R1072 vdd vdd 0.001
R1073 vdd vdd 0.001
R108 A:F171 A:F335 1643.25
R109 A:F171 A:F331 8699.01
R11 vdd vdd 0.001
R110 A:F171 A:F183 6439.37
R111 A:F171 A:F179 1845.53
R112 A:F171 A:F175 563.846
R113 A:F171 A:F3 162.829
R114 A:F175 A:F355 1375.65
R115 A:F175 A:F351 381.063
R116 A:F175 A:F347 115.236
R117 A:F175 A:F343 490.301
R118 A:F175 A:F339 2069.79
R119 A:F175 A:F335 5641.18
R12 vdd vdd 0.001
R120 A:F175 A:F183 1582
R121 A:F175 A:F179 438.223
R122 A:F175 A:F3 137.153
R123 A:F179 A:F355 373.944
R124 A:F179 A:F351 100.972
R125 A:F179 A:F347 377.773
R126 A:F179 A:F343 1604.81
R127 A:F179 A:F339 6774.68
R128 A:F179 A:F183 430.036
R129 A:F179 A:F3 204.153
R13 vdd vdd 0.001
R130 A:F323 A:F339 21379.6
R131 A:F323 A:F335 6762.83
R132 A:F323 A:F331 1276.78
R133 A:F323 A:F327 352.733
R134 A:F323 A:F319 361.284
R135 A:F323 A:F315 1038.84
R136 A:F323 A:F155 405.643
R137 A:F323 A:F147 361.284
R138 A:F323 A:F143 1038.84
R139 A:F323 A:F3 1589.08
R14 vdd vdd 0.001
R140 A:F327 A:F343 10480
R141 A:F327 A:F339 4315.85
R142 A:F327 A:F335 1523.83
R143 A:F327 A:F331 308.828
R144 A:F327 A:F319 1245.32
R145 A:F327 A:F315 3580.81
R146 A:F327 A:F155 98.1172
R147 A:F327 A:F147 1245.32
R148 A:F327 A:F143 3580.81
R149 A:F327 A:F3 384.367
R15 vdd vdd 0.001
R150 A:F331 A:F343 7477.04
R151 A:F331 A:F339 1655.9
R152 A:F331 A:F335 523.797
R153 A:F331 A:F319 4507.64
R154 A:F331 A:F315 12961.3
R155 A:F331 A:F155 355.152
R156 A:F331 A:F147 4507.64
R157 A:F331 A:F143 12961.3
R158 A:F331 A:F3 124.007
R159 A:F315 A:F319 286.499
R16 vdd vdd 0.001
R160 A:F315 A:F155 4117.93
R161 A:F315 A:F147 286.499
R162 A:F315 A:F143 79.5284
R163 A:F315 A:F3 16131.7
R164 A:F335 A:F347 6628.86
R165 A:F335 A:F343 1428.32
R166 A:F335 A:F339 330.367
R167 A:F335 A:F155 1867.97
R168 A:F335 A:F147 13114
R169 A:F335 A:F3 113.375
R17 vdd vdd 0.001
R170 A:F319 A:F155 1432.11
R171 A:F319 A:F147 99.6374
R172 A:F319 A:F143 286.499
R173 A:F319 A:F3 5610.21
R174 A:F339 A:F355 20554.8
R175 A:F339 A:F351 5891.02
R176 A:F339 A:F347 1799.82
R177 A:F339 A:F343 387.955
R178 A:F339 A:F155 5905.29
R179 A:F339 A:F3 175.733
R18 vdd vdd 0.001
R180 A:F343 A:F355 4869.09
R181 A:F343 A:F351 1395.49
R182 A:F343 A:F347 426.348
R183 A:F343 A:F183 5599.45
R184 A:F343 A:F155 14339.5
R185 A:F343 A:F3 141.566
R186 A:F155 A:F147 1432.11
R187 A:F155 A:F143 4117.93
R188 A:F155 A:F3 442.023
R189 A:F347 A:F355 1101.35
R19 vdd vdd 0.001
R190 A:F347 A:F351 328.498
R191 A:F347 A:F183 1266.55
R192 A:F347 A:F3 119.264
R193 A:F351 A:F355 325.169
R194 A:F351 A:F183 373.944
R195 A:F351 A:F3 177.525
R196 A:F355 A:F183 82.0527
R197 A:F355 A:F3 167.405
R198 A:F183 A:F3 190.961
R199 A:F3 A:F147 5610.21
R2 vdd vdd 0.001
R20 vdd vdd 0.001
R200 A:F3 A:F143 16131.7
R201 A:F143 A:F147 286.499
R202 gnd gnd 0.001
R203 gnd gnd 0.001
R204 gnd gnd 0.001
R205 gnd gnd 0.001
R206 gnd gnd 0.001
R207 gnd gnd 0.001
R208 gnd gnd 0.001
R209 gnd gnd 0.001
R21 vdd vdd 0.001
R210 gnd gnd 0.001
R211 gnd gnd 0.001
R212 gnd gnd 0.001
R213 gnd gnd 0.001
R214 gnd gnd 0.001
R215 gnd gnd 0.001
R216 gnd gnd 0.001
R217 gnd gnd 0.001
R218 gnd gnd 0.001
R219 gnd gnd 0.001
R22 vdd vdd 0.001
R220 gnd gnd 0.001
R221 gnd gnd 0.001
R222 gnd gnd 0.001
R223 gnd gnd 0.001
R224 gnd gnd 0.001
R225 gnd gnd 0.001
R226 gnd gnd 0.001
R227 gnd gnd 0.001
R228 gnd gnd 0.001
R229 gnd gnd 0.001
R23 vdd vdd 0.001
R230 gnd gnd 0.001
R231 gnd gnd 0.001
R232 gnd gnd 0.001
R233 gnd gnd 0.001
R234 gnd gnd 0.001
R235 gnd gnd 0.001
R236 gnd gnd 0.001
R237 gnd gnd 0.001
R238 gnd gnd 0.001
R239 gnd gnd 0.001
R24 vdd vdd 0.001
R240 gnd gnd 0.001
R241 gnd gnd 0.001
R242 gnd gnd 0.001
R243 gnd gnd 0.001
R244 gnd gnd 0.001
R245 gnd gnd 0.001
R246 gnd gnd 0.0256454
R247 gnd gnd 37.6237
R248 Z Z:F4 0.001
R249 Z:F4 Z:F266 94.9766
R25 vdd vdd 0.001
R250 Z:F4 Z:F258 51.4203
R251 Z:F4 Z:F256 35.2747
R252 Z:F4 Z:F248 26.5644
R253 Z:F4 Z:F240 18.822
R254 Z:F4 Z:F232 18.8025
R255 Z:F4 Z:F224 25.7475
R256 Z:F4 Z:F216 34.7326
R257 Z:F4 Z:F208 52.5367
R258 Z:F4 Z:F200 105.603
R259 Z:F4 Z:F94 94.3663
R26 vdd vdd 0.001
R260 Z:F4 Z:F86 51.3507
R261 Z:F4 Z:F78 35.4039
R262 Z:F4 Z:F70 26.5449
R263 Z:F4 Z:F62 18.8547
R264 Z:F4 Z:F54 18.8449
R265 Z:F4 Z:F46 25.8417
R266 Z:F4 Z:F38 34.802
R267 Z:F4 Z:F30 52.729
R268 Z:F4 Z:F22 105.99
R269 Z:F4 Z:148 0.533397
R27 vdd vdd 0.001
R270 Z:F4 Z:1616 0.58015
R271 Z:F258 Z:F264 0.001
R272 Z:F258 Z:1616 30.4599
R273 Z:F306 Z:F312 0.001
R274 Z:F306 Z:F298 644.033
R275 Z:F306 Z:F296 1020.85
R276 Z:F306 Z:F282 2393.77
R277 Z:F306 Z:1616 20.7299
R278 Z:1616 Z:F298 20.4933
R279 Z:1616 Z:F296 20.0333
R28 vdd vdd 0.001
R280 Z:1616 Z:F282 19.3127
R281 Z:1616 Z:F274 18.7825
R282 Z:1616 Z:F266 23.7242
R283 Z:1616 Z:F256 43.5412
R284 Z:1616 Z:F248 67.1123
R285 Z:1616 Z:F134 22.1366
R286 Z:1616 Z:F126 21.7176
R287 Z:1616 Z:F124 20.9181
R288 Z:1616 Z:F110 19.7
R289 Z:1616 Z:F102 18.8027
R29 vdd vdd 0.001
R290 Z:1616 Z:F94 23.7881
R291 Z:1616 Z:F86 30.6614
R292 Z:1616 Z:F78 42.9936
R293 Z:1616 Z:F70 66.7189
R294 Z:148 Z:F224 76.0559
R295 Z:148 Z:F216 42.4658
R296 Z:148 Z:F208 30.261
R297 Z:148 Z:F200 23.0589
R298 Z:148 Z:F192 18.75
R299 Z:148 Z:F46 74.7851
R3 vdd vdd 0.001
R30 vdd vdd 0.001
R300 Z:148 Z:F38 42.4369
R301 Z:148 Z:F30 30.0708
R302 Z:148 Z:F22 22.994
R303 Z:148 Z:F14 18.8187
R304 Z:F134 Z:F140 0.001
R305 Z:F134 Z:F126 407.901
R306 Z:F134 Z:F124 650.29
R307 Z:F134 Z:F110 1529.89
R308 Z:F266 Z:F272 0.001
R309 Z:F274 Z:F280 0.001
R31 vdd vdd 0.001
R310 Z:F232 Z:F226 0.001
R311 Z:F54 Z:F60 0.001
R312 Z:F192 Z:F186 0.001
R313 Z:F240 Z:F234 0.001
R314 Z:F248 Z:F242 0.001
R315 Z:F256 Z:F250 0.001
R316 Z:F282 Z:F298 2366.44
R317 Z:F282 Z:F296 3751.01
R318 Z:F282 Z:F288 0.001
R319 Z:F296 Z:F298 1009.2
R32 vdd vdd 0.001
R320 Z:F296 Z:F290 0.001
R321 Z:F298 Z:F304 0.001
R322 Z:F14 Z:F20 0.001
R323 Z:F62 Z:F68 0.001
R324 Z:F70 Z:F76 0.001
R325 Z:F78 Z:F84 0.001
R326 Z:F86 Z:F92 0.001
R327 Z:F94 Z:F100 0.001
R328 Z:F102 Z:F108 0.001
R329 Z:F110 Z:F126 1500.93
R33 vdd vdd 0.001
R330 Z:F110 Z:F124 2392.84
R331 Z:F110 Z:F116 0.001
R332 Z:F124 Z:F126 637.981
R333 Z:F124 Z:F118 0.001
R334 Z:F126 Z:F132 0.001
R335 Z:F200 Z:F194 0.001
R336 Z:F208 Z:F202 0.001
R337 Z:F216 Z:F210 0.001
R338 Z:F224 Z:F218 0.001
R339 Z:F22 Z:F28 0.001
R34 vdd vdd 0.001
R340 Z:F30 Z:F36 0.001
R341 Z:F38 Z:F44 0.001
R342 Z:F46 Z:F52 0.001
R343 gnd gnd 0.001
R344 gnd gnd 61.2192
R345 gnd gnd 28.7826
R346 gnd gnd 18.8094
R347 gnd gnd 21.0316
R348 gnd gnd 23.6222
R349 gnd gnd 26.8547
R35 vdd vdd 0.001
R350 gnd gnd 30.7922
R351 gnd gnd 35.7333
R352 gnd gnd 42.4131
R353 gnd gnd 51.1125
R354 gnd gnd 64.4914
R355 gnd gnd 87.9549
R356 gnd gnd 129.147
R357 gnd gnd 259.276
R358 gnd gnd 1.76874
R359 gnd gnd 0.370054
R36 vdd vdd 0.001
R360 gnd gnd 4.05225
R361 gnd gnd 7.84885
R362 gnd gnd 13.3537
R363 gnd gnd 233.94
R364 gnd gnd 122.449
R365 gnd gnd 86.8148
R366 gnd gnd 58.9481
R367 gnd gnd 51.031
R368 gnd gnd 42.1248
R369 gnd gnd 34.664
R37 vdd vdd 0.001
R370 gnd gnd 30.116
R371 gnd gnd 26.7231
R372 gnd gnd 23.1385
R373 gnd gnd 20.4097
R374 gnd gnd 18.8269
R375 gnd gnd 0.001
R376 gnd gnd 18.8134
R377 gnd gnd 2337.13
R378 gnd gnd 3902.68
R379 gnd gnd 3859.44
R38 vdd vdd 0.001
R380 gnd gnd 3796.06
R381 gnd gnd 0.001
R382 gnd gnd 19.3478
R383 gnd gnd 1922.39
R384 gnd gnd 1911.41
R385 gnd gnd 1890.23
R386 gnd gnd 1859.18
R387 gnd gnd 0.001
R388 gnd gnd 19.9047
R389 gnd gnd 1263.24
R39 vdd vdd 0.001
R390 gnd gnd 1256.02
R391 gnd gnd 1242.1
R392 gnd gnd 0.001
R393 gnd gnd 20.3434
R394 gnd gnd 1284.33
R395 gnd gnd 733.939
R396 gnd gnd 0.001
R397 gnd gnd 20.6831
R398 gnd gnd 741.086
R399 gnd gnd 0.001
R4 vdd vdd 0.001
R40 vdd vdd 0.001
R400 gnd gnd 20.9148
R401 gnd gnd 0.001
R402 gnd gnd 21.035
R403 gnd gnd 27.3976
R404 gnd gnd 54.9796
R405 gnd gnd 1340.05
R406 gnd gnd 1223.85
R407 gnd gnd 0.001
R408 gnd gnd 1111.97
R409 gnd gnd 659.944
R41 vdd vdd 0.001
R410 gnd gnd 0.001
R411 gnd gnd 670.539
R412 gnd gnd 673.866
R413 gnd gnd 805.257
R414 gnd gnd 1333.65
R415 gnd gnd 936.842
R416 gnd gnd 0.001
R417 gnd gnd 1220.45
R418 gnd gnd 0.001
R419 gnd gnd 1382.98
R42 vdd vdd 0.001
R420 gnd gnd 0.001
R421 gnd gnd 1312.65
R422 gnd gnd 0.001
R423 gnd gnd 0.001
R424 gnd gnd 0.001
R425 gnd gnd 0.001
R426 gnd gnd 0.001
R427 gnd gnd 0.001
R428 gnd gnd 0.001
R429 gnd gnd 0.001
R43 vdd vdd 0.001
R430 gnd gnd 0.001
R431 net0513:1020 net0513:F354 39.4881
R432 net0513:1020 net0513:F346 38.363
R433 net0513:1020 net0513:F338 36.3666
R434 net0513:1020 net0513:F330 33.6764
R435 net0513:1020 net0513:F322 30.261
R436 net0513:1020 net0513:F314 27.2833
R437 net0513:1020 net0513:F311 466.551
R438 net0513:1020 net0513:F307 150.29
R439 net0513:1020 net0513:F303 273.995
R44 vdd vdd 0.001
R440 net0513:1020 net0513:F299 159.147
R441 net0513:1020 net0513:F295 1000.2
R442 net0513:1020 net0513:F291 706.045
R443 net0513:1020 net0513:F287 174.365
R444 net0513:1020 net0513:F283 653.06
R445 net0513:1020 net0513:F279 2315.84
R446 net0513:1020 net0513:F275 8820.33
R447 net0513:1020 net0513:F182 39.8273
R448 net0513:1020 net0513:F174 38.6296
R449 net0513:1020 net0513:F166 36.5053
R45 vdd vdd 37.6252
R450 net0513:1020 net0513:F158 33.6845
R451 net0513:1020 net0513:F150 29.9597
R452 net0513:1020 net0513:F142 26.7791
R453 net0513:1020 net0513:F139 466.551
R454 net0513:1020 net0513:F135 150.29
R455 net0513:1020 net0513:F131 273.995
R456 net0513:1020 net0513:F127 159.147
R457 net0513:1020 net0513:F123 1000.2
R458 net0513:1020 net0513:F119 706.045
R459 net0513:1020 net0513:F115 174.365
R46 A A:F3 0.001
R460 net0513:1020 net0513:F111 653.06
R461 net0513:1020 net0513:F107 2315.84
R462 net0513:1020 net0513:F103 8820.33
R463 net0513:1020 net0513:744 7976.65
R464 net0513:1020 net0513:924 32.2937
R465 net0513:924 net0513:F311 9208.95
R466 net0513:924 net0513:F307 2966.47
R467 net0513:924 net0513:F303 828.521
R468 net0513:924 net0513:F299 248.324
R469 net0513:924 net0513:F295 53.6837
R47 A:F151 A:F343 25957.5
R470 net0513:924 net0513:F291 77.832
R471 net0513:924 net0513:F287 291.382
R472 net0513:924 net0513:F283 1091.33
R473 net0513:924 net0513:F279 3870
R474 net0513:924 net0513:F275 14739.7
R475 net0513:924 net0513:F139 9208.95
R476 net0513:924 net0513:F135 2966.47
R477 net0513:924 net0513:F131 828.521
R478 net0513:924 net0513:F127 248.324
R479 net0513:924 net0513:F123 53.6837
R48 A:F151 A:F339 21379.6
R480 net0513:924 net0513:F119 77.832
R481 net0513:924 net0513:F115 291.382
R482 net0513:924 net0513:F111 1091.33
R483 net0513:924 net0513:F107 3870
R484 net0513:924 net0513:F103 14739.7
R485 net0513:924 net0513:744 13329.8
R486 net0513:744 net0513:F291 23429.3
R487 net0513:744 net0513:F287 5786.11
R488 net0513:744 net0513:F283 1260.64
R489 net0513:744 net0513:F279 357.269
R49 A:F151 A:F335 6762.83
R490 net0513:744 net0513:F275 101.345
R491 net0513:744 net0513:F271 28.75
R492 net0513:744 net0513:F267 101.341
R493 net0513:744 net0513:F263 357.105
R494 net0513:744 net0513:F259 1258.76
R495 net0513:744 net0513:F255 4435.61
R496 net0513:744 net0513:F251 15635.1
R497 net0513:744 net0513:F119 23429.3
R498 net0513:744 net0513:F115 5786.11
R499 net0513:744 net0513:F111 1260.64
R5 vdd vdd 0.001
R50 A:F151 A:F331 1276.78
R500 net0513:744 net0513:F107 357.269
R501 net0513:744 net0513:F103 101.345
R502 net0513:744 net0513:F99 28.75
R503 net0513:744 net0513:F95 101.341
R504 net0513:744 net0513:F91 357.105
R505 net0513:744 net0513:F87 1258.76
R506 net0513:744 net0513:F83 4435.61
R507 net0513:744 net0513:F79 15635.1
R508 net0513:F303 net0513:F311 1241.93
R509 net0513:F303 net0513:F307 400.061
R51 A:F151 A:F327 352.733
R510 net0513:F303 net0513:F299 427.964
R511 net0513:F303 net0513:F295 2689.66
R512 net0513:F303 net0513:F139 1241.93
R513 net0513:F303 net0513:F135 400.061
R514 net0513:F303 net0513:F131 111.735
R515 net0513:F303 net0513:F127 427.964
R516 net0513:F303 net0513:F123 2689.66
R517 net0513:F307 net0513:F311 385.755
R518 net0513:F307 net0513:F299 1532.3
R519 net0513:F307 net0513:F295 9630.15
R52 A:F151 A:F323 102.333
R520 net0513:F307 net0513:F139 385.755
R521 net0513:F307 net0513:F135 124.263
R522 net0513:F307 net0513:F131 400.061
R523 net0513:F307 net0513:F127 1532.3
R524 net0513:F307 net0513:F123 9630.15
R525 net0513:F311 net0513:F299 4756.78
R526 net0513:F311 net0513:F139 79.2134
R527 net0513:F311 net0513:F135 385.755
R528 net0513:F311 net0513:F131 1241.93
R529 net0513:F311 net0513:F127 4756.78
R53 A:F151 A:F319 361.284
R530 net0513:F314 net0513:F354 646.763
R531 net0513:F314 net0513:F346 628.335
R532 net0513:F314 net0513:F338 595.636
R533 net0513:F314 net0513:F330 551.574
R534 net0513:F314 net0513:F322 495.635
R535 net0513:F314 net0513:F320 0.001
R536 net0513:F314 net0513:F182 1254.94
R537 net0513:F314 net0513:F174 1217.2
R538 net0513:F314 net0513:F166 1150.27
R539 net0513:F314 net0513:F158 1061.39
R54 A:F151 A:F315 1038.84
R540 net0513:F314 net0513:F150 958.854
R541 net0513:F314 net0513:F142 843.799
R542 net0513:F295 net0513:F299 806.144
R543 net0513:F295 net0513:F139 14947.7
R544 net0513:F295 net0513:F135 9630.15
R545 net0513:F295 net0513:F131 2689.66
R546 net0513:F295 net0513:F127 806.144
R547 net0513:F295 net0513:F123 171.584
R548 net0513:F79 net0513:F267 17288.8
R549 net0513:F79 net0513:F263 4539.31
R55 A:F151 A:F167 24183.1
R550 net0513:F79 net0513:F259 1280.51
R551 net0513:F79 net0513:F255 363.1
R552 net0513:F79 net0513:F251 103.038
R553 net0513:F79 net0513:F247 363.085
R554 net0513:F79 net0513:F243 1279.84
R555 net0513:F79 net0513:F239 3930.08
R556 net0513:F79 net0513:F235 13853.6
R557 net0513:F79 net0513:F95 17288.8
R558 net0513:F79 net0513:F91 4539.31
R559 net0513:F79 net0513:F87 1280.51
R56 A:F151 A:F163 7786.31
R560 net0513:F79 net0513:F83 363.1
R561 net0513:F79 net0513:F75 363.085
R562 net0513:F79 net0513:F71 1279.84
R563 net0513:F79 net0513:F67 3930.08
R564 net0513:F79 net0513:F63 13853.6
R565 net0513:F103 net0513:F291 12953.7
R566 net0513:F103 net0513:F287 6398.11
R567 net0513:F103 net0513:F283 1393.97
R568 net0513:F103 net0513:F279 395.057
R569 net0513:F103 net0513:F275 112.064
R57 A:F151 A:F159 1468.29
R570 net0513:F103 net0513:F119 12953.7
R571 net0513:F103 net0513:F115 6398.11
R572 net0513:F103 net0513:F111 1393.97
R573 net0513:F103 net0513:F107 395.057
R574 net0513:F191 net0513:F207 12305.1
R575 net0513:F191 net0513:F203 4477.44
R576 net0513:F191 net0513:F199 1269.58
R577 net0513:F191 net0513:F195 360.151
R578 net0513:F191 net0513:F187 276.803
R579 net0513:F191 net0513:F35 15877.6
R58 A:F151 A:F155 405.643
R580 net0513:F191 net0513:F31 3899.93
R581 net0513:F191 net0513:F27 1269.58
R582 net0513:F191 net0513:F23 360.151
R583 net0513:F191 net0513:F19 95.9508
R584 net0513:F191 net0513:F15 265.731
R585 net0513:F299 net0513:F139 4756.78
R586 net0513:F299 net0513:F135 1532.3
R587 net0513:F299 net0513:F131 427.964
R588 net0513:F299 net0513:F127 128.269
R589 net0513:F299 net0513:F123 806.144
R59 A:F151 A:F147 361.284
R590 net0513:F83 net0513:F267 4904.76
R591 net0513:F83 net0513:F263 1287.78
R592 net0513:F83 net0513:F259 363.274
R593 net0513:F83 net0513:F255 103.01
R594 net0513:F83 net0513:F251 363.1
R595 net0513:F83 net0513:F247 1279.49
R596 net0513:F83 net0513:F243 4510.07
R597 net0513:F83 net0513:F239 15995.6
R598 net0513:F83 net0513:F235 24618.6
R599 net0513:F83 net0513:F95 4904.76
R6 vdd vdd 0.001
R60 A:F151 A:F143 1038.84
R600 net0513:F83 net0513:F91 1287.78
R601 net0513:F83 net0513:F87 363.274
R602 net0513:F83 net0513:F75 1279.49
R603 net0513:F83 net0513:F71 4510.07
R604 net0513:F83 net0513:F67 15995.6
R605 net0513:F83 net0513:F63 24618.6
R606 net0513:F107 net0513:F291 6802.18
R607 net0513:F107 net0513:F287 1679.87
R608 net0513:F107 net0513:F283 365.997
R609 net0513:F107 net0513:F279 103.725
R61 A:F151 A:F3 1589.08
R610 net0513:F107 net0513:F275 395.057
R611 net0513:F107 net0513:F119 6802.18
R612 net0513:F107 net0513:F115 1679.87
R613 net0513:F107 net0513:F111 365.997
R614 net0513:F199 net0513:F215 15905.4
R615 net0513:F199 net0513:F211 4513.67
R616 net0513:F199 net0513:F207 1280.5
R617 net0513:F199 net0513:F203 363.264
R618 net0513:F199 net0513:F195 363.623
R619 net0513:F199 net0513:F187 3516.04
R62 A:F159 A:F343 8598.59
R620 net0513:F199 net0513:F43 15905.4
R621 net0513:F199 net0513:F39 3887.96
R622 net0513:F199 net0513:F35 1261.9
R623 net0513:F199 net0513:F31 362.916
R624 net0513:F199 net0513:F27 103.053
R625 net0513:F199 net0513:F23 363.623
R626 net0513:F199 net0513:F19 1218.8
R627 net0513:F199 net0513:F15 3375.4
R628 net0513:F322 net0513:F354 413.662
R629 net0513:F322 net0513:F346 401.876
R63 A:F159 A:F339 1904.28
R630 net0513:F322 net0513:F338 380.962
R631 net0513:F322 net0513:F330 423.966
R632 net0513:F322 net0513:F328 0.001
R633 net0513:F322 net0513:F182 1391.91
R634 net0513:F322 net0513:F174 1350.05
R635 net0513:F322 net0513:F166 1275.81
R636 net0513:F322 net0513:F158 1177.22
R637 net0513:F322 net0513:F150 1063.5
R638 net0513:F322 net0513:F142 935.891
R639 net0513:F127 net0513:F139 4756.78
R64 A:F159 A:F335 602.366
R640 net0513:F127 net0513:F135 1532.3
R641 net0513:F127 net0513:F131 427.964
R642 net0513:F127 net0513:F123 806.144
R643 net0513:F87 net0513:F267 1391.9
R644 net0513:F87 net0513:F263 365.453
R645 net0513:F87 net0513:F259 103.092
R646 net0513:F87 net0513:F255 363.274
R647 net0513:F87 net0513:F251 1280.51
R648 net0513:F87 net0513:F247 3930.07
R649 net0513:F87 net0513:F243 13853.1
R65 A:F159 A:F331 114.581
R650 net0513:F87 net0513:F95 1391.9
R651 net0513:F87 net0513:F91 365.453
R652 net0513:F87 net0513:F75 3930.07
R653 net0513:F87 net0513:F71 13853.1
R654 net0513:F111 net0513:F291 1918.19
R655 net0513:F111 net0513:F287 473.717
R656 net0513:F111 net0513:F283 103.21
R657 net0513:F111 net0513:F279 365.997
R658 net0513:F111 net0513:F275 1393.97
R659 net0513:F111 net0513:F119 1918.19
R66 A:F159 A:F327 355.152
R660 net0513:F111 net0513:F115 473.717
R661 net0513:F207 net0513:F223 16007
R662 net0513:F207 net0513:F219 4513.92
R663 net0513:F207 net0513:F215 1279.93
R664 net0513:F207 net0513:F211 363.222
R665 net0513:F207 net0513:F203 363.234
R666 net0513:F207 net0513:F195 4518.26
R667 net0513:F207 net0513:F51 16007
R668 net0513:F207 net0513:F47 4513.92
R669 net0513:F207 net0513:F43 1279.93
R67 A:F159 A:F323 1468.29
R670 net0513:F207 net0513:F39 363.222
R671 net0513:F207 net0513:F35 103.044
R672 net0513:F207 net0513:F31 363.234
R673 net0513:F207 net0513:F27 1280.5
R674 net0513:F207 net0513:F23 4518.26
R675 net0513:F207 net0513:F19 11812.9
R676 net0513:F330 net0513:F354 300.484
R677 net0513:F330 net0513:F346 291.922
R678 net0513:F330 net0513:F338 276.731
R679 net0513:F330 net0513:F336 0.001
R68 A:F159 A:F319 5183.79
R680 net0513:F330 net0513:F182 1549
R681 net0513:F330 net0513:F174 1502.42
R682 net0513:F330 net0513:F166 1419.8
R683 net0513:F330 net0513:F158 1310.09
R684 net0513:F330 net0513:F150 1183.53
R685 net0513:F330 net0513:F142 1041.52
R686 net0513:F338 net0513:F354 230.15
R687 net0513:F338 net0513:F346 223.592
R688 net0513:F338 net0513:F344 0.001
R689 net0513:F338 net0513:F182 1672.74
R69 A:F159 A:F315 14905.6
R690 net0513:F338 net0513:F174 1622.44
R691 net0513:F338 net0513:F166 1533.22
R692 net0513:F338 net0513:F158 1414.75
R693 net0513:F338 net0513:F150 1278.08
R694 net0513:F338 net0513:F142 1124.72
R695 net0513:F346 net0513:F354 182.381
R696 net0513:F346 net0513:F352 0.001
R697 net0513:F346 net0513:F182 1764.57
R698 net0513:F346 net0513:F174 1711.51
R699 net0513:F346 net0513:F166 1617.39
R7 vdd vdd 0.001
R70 A:F159 A:F171 10003.9
R700 net0513:F346 net0513:F158 1492.41
R701 net0513:F346 net0513:F150 1348.24
R702 net0513:F346 net0513:F142 1186.46
R703 net0513:F354 net0513:F182 1816.32
R704 net0513:F354 net0513:F174 1761.7
R705 net0513:F354 net0513:F166 1664.82
R706 net0513:F354 net0513:F158 1536.18
R707 net0513:F354 net0513:F150 1387.78
R708 net0513:F354 net0513:F142 1221.26
R709 net0513:F131 net0513:F139 1241.93
R71 A:F159 A:F167 2153.99
R710 net0513:F131 net0513:F135 400.061
R711 net0513:F131 net0513:F123 2689.66
R712 net0513:F135 net0513:F139 385.755
R713 net0513:F135 net0513:F123 9630.15
R714 net0513:F91 net0513:F267 394.875
R715 net0513:F91 net0513:F263 103.677
R716 net0513:F91 net0513:F259 365.453
R717 net0513:F91 net0513:F255 1287.78
R718 net0513:F91 net0513:F251 4539.31
R719 net0513:F91 net0513:F247 15995.5
R72 A:F159 A:F163 693.528
R720 net0513:F91 net0513:F243 24617.8
R721 net0513:F91 net0513:F95 394.875
R722 net0513:F91 net0513:F75 15995.5
R723 net0513:F91 net0513:F71 24617.8
R724 net0513:F95 net0513:F267 112.06
R725 net0513:F95 net0513:F263 394.875
R726 net0513:F95 net0513:F259 1391.9
R727 net0513:F95 net0513:F255 4904.76
R728 net0513:F95 net0513:F251 17288.8
R729 net0513:F115 net0513:F291 512.152
R73 A:F159 A:F155 408.425
R730 net0513:F115 net0513:F287 126.481
R731 net0513:F115 net0513:F283 473.717
R732 net0513:F115 net0513:F279 1679.87
R733 net0513:F115 net0513:F275 6398.11
R734 net0513:F115 net0513:F119 512.152
R735 net0513:F119 net0513:F291 131.957
R736 net0513:F119 net0513:F287 512.152
R737 net0513:F119 net0513:F283 1918.19
R738 net0513:F119 net0513:F279 6802.18
R739 net0513:F279 net0513:F291 6802.18
R74 A:F159 A:F147 5183.79
R740 net0513:F279 net0513:F287 1679.87
R741 net0513:F279 net0513:F283 365.997
R742 net0513:F279 net0513:F275 395.057
R743 net0513:F287 net0513:F291 512.152
R744 net0513:F287 net0513:F283 473.717
R745 net0513:F287 net0513:F275 6398.11
R746 net0513:F275 net0513:F283 1393.97
R747 net0513:F139 net0513:F123 14947.7
R748 net0513:F215 net0513:F231 12405.8
R749 net0513:F215 net0513:F227 4513.59
R75 A:F159 A:F143 14905.6
R750 net0513:F215 net0513:F223 1279.93
R751 net0513:F215 net0513:F219 363.077
R752 net0513:F215 net0513:F211 363.084
R753 net0513:F215 net0513:F203 4511.79
R754 net0513:F215 net0513:F59 16007.6
R755 net0513:F215 net0513:F55 3931.48
R756 net0513:F215 net0513:F51 1279.93
R757 net0513:F215 net0513:F47 363.085
R758 net0513:F215 net0513:F43 103.002
R759 net0513:F215 net0513:F39 363.084
R76 A:F159 A:F3 142.608
R760 net0513:F215 net0513:F35 1279.93
R761 net0513:F215 net0513:F31 4511.79
R762 net0513:F215 net0513:F27 15905.4
R763 net0513:F219 net0513:F235 15222.4
R764 net0513:F219 net0513:F231 4316.44
R765 net0513:F219 net0513:F227 1224.34
R766 net0513:F219 net0513:F223 363.113
R767 net0513:F219 net0513:F211 1279.85
R768 net0513:F219 net0513:F203 15911.7
R769 net0513:F219 net0513:F67 23560.9
R77 A:F163 A:F347 7623.19
R770 net0513:F219 net0513:F63 13258.4
R771 net0513:F219 net0513:F59 4316.44
R772 net0513:F219 net0513:F55 1224.34
R773 net0513:F219 net0513:F51 363.113
R774 net0513:F219 net0513:F47 103.039
R775 net0513:F219 net0513:F43 363.077
R776 net0513:F219 net0513:F39 1279.85
R777 net0513:F219 net0513:F35 4513.92
R778 net0513:F219 net0513:F31 15911.7
R779 net0513:F223 net0513:F239 12406.2
R78 A:F163 A:F343 1642.56
R780 net0513:F223 net0513:F235 4515.78
R781 net0513:F223 net0513:F231 1280.49
R782 net0513:F223 net0513:F227 363.206
R783 net0513:F223 net0513:F211 4511.76
R784 net0513:F223 net0513:F67 16008.1
R785 net0513:F223 net0513:F63 3933.16
R786 net0513:F223 net0513:F59 1280.49
R787 net0513:F223 net0513:F55 363.206
R788 net0513:F223 net0513:F51 103.044
R789 net0513:F223 net0513:F47 363.22
R79 A:F163 A:F339 379.922
R790 net0513:F223 net0513:F43 1279.93
R791 net0513:F223 net0513:F39 4511.76
R792 net0513:F223 net0513:F35 16007
R793 net0513:F227 net0513:F243 15897.3
R794 net0513:F227 net0513:F239 4507.81
R795 net0513:F227 net0513:F235 1279.2
R796 net0513:F227 net0513:F231 362.902
R797 net0513:F227 net0513:F211 15910.5
R798 net0513:F227 net0513:F75 24605.5
R799 net0513:F227 net0513:F71 13846.2
R8 vdd vdd 0.001
R80 A:F163 A:F335 114.473
R800 net0513:F227 net0513:F67 4507.81
R801 net0513:F227 net0513:F63 1279.2
R802 net0513:F227 net0513:F59 362.902
R803 net0513:F227 net0513:F55 103.029
R804 net0513:F227 net0513:F51 363.206
R805 net0513:F227 net0513:F47 1280.27
R806 net0513:F227 net0513:F43 4513.59
R807 net0513:F227 net0513:F39 15910.5
R808 net0513:F231 net0513:F247 12401.6
R809 net0513:F231 net0513:F243 4514.11
R81 A:F163 A:F331 603.067
R810 net0513:F231 net0513:F239 1280.02
R811 net0513:F231 net0513:F235 363.236
R812 net0513:F231 net0513:F75 16002.2
R813 net0513:F231 net0513:F71 3931.7
R814 net0513:F231 net0513:F67 1280.02
R815 net0513:F231 net0513:F63 363.236
R816 net0513:F231 net0513:F59 103.048
R817 net0513:F231 net0513:F55 362.902
R818 net0513:F231 net0513:F51 1280.49
R819 net0513:F231 net0513:F47 4513.6
R82 A:F163 A:F327 1754.45
R820 net0513:F231 net0513:F43 12405.8
R821 net0513:F235 net0513:F251 15905.8
R822 net0513:F235 net0513:F247 4510.22
R823 net0513:F235 net0513:F243 1279.89
R824 net0513:F235 net0513:F239 363.097
R825 net0513:F235 net0513:F75 4510.22
R826 net0513:F235 net0513:F71 1279.89
R827 net0513:F235 net0513:F67 363.097
R828 net0513:F235 net0513:F63 103.042
R829 net0513:F235 net0513:F59 363.236
R83 A:F163 A:F323 7786.31
R830 net0513:F235 net0513:F55 1279.2
R831 net0513:F235 net0513:F51 4515.78
R832 net0513:F235 net0513:F47 15917.7
R833 net0513:F239 net0513:F255 12396.5
R834 net0513:F239 net0513:F251 4512.25
R835 net0513:F239 net0513:F247 1279.49
R836 net0513:F239 net0513:F243 363.087
R837 net0513:F239 net0513:F75 1279.49
R838 net0513:F239 net0513:F71 363.087
R839 net0513:F239 net0513:F67 103.006
R84 A:F163 A:F175 6487.36
R840 net0513:F239 net0513:F63 363.097
R841 net0513:F239 net0513:F59 1280.02
R842 net0513:F239 net0513:F55 4507.81
R843 net0513:F239 net0513:F51 12406.2
R844 net0513:F243 net0513:F259 15905.2
R845 net0513:F243 net0513:F255 4510.07
R846 net0513:F243 net0513:F251 1279.84
R847 net0513:F243 net0513:F247 363.084
R848 net0513:F243 net0513:F75 363.084
R849 net0513:F243 net0513:F71 103.038
R85 A:F163 A:F171 1889.74
R850 net0513:F243 net0513:F67 363.087
R851 net0513:F243 net0513:F63 1279.89
R852 net0513:F243 net0513:F59 4514.11
R853 net0513:F243 net0513:F55 15897.3
R854 net0513:F247 net0513:F263 12396.5
R855 net0513:F247 net0513:F259 4512.23
R856 net0513:F247 net0513:F255 1279.49
R857 net0513:F247 net0513:F251 363.085
R858 net0513:F247 net0513:F75 103.005
R859 net0513:F247 net0513:F71 363.084
R86 A:F163 A:F167 436.909
R860 net0513:F247 net0513:F67 1279.49
R861 net0513:F247 net0513:F63 4510.22
R862 net0513:F247 net0513:F59 12401.6
R863 net0513:F255 net0513:F267 4904.76
R864 net0513:F255 net0513:F263 1287.78
R865 net0513:F255 net0513:F259 363.274
R866 net0513:F255 net0513:F251 363.1
R867 net0513:F255 net0513:F75 1279.49
R868 net0513:F255 net0513:F71 4510.07
R869 net0513:F255 net0513:F67 12396.5
R87 A:F163 A:F155 2150.67
R870 net0513:F263 net0513:F267 394.875
R871 net0513:F263 net0513:F259 365.453
R872 net0513:F263 net0513:F251 4539.31
R873 net0513:F263 net0513:F75 12396.5
R874 net0513:F259 net0513:F267 1391.9
R875 net0513:F259 net0513:F251 1280.51
R876 net0513:F259 net0513:F75 4512.23
R877 net0513:F259 net0513:F71 15905.2
R878 net0513:F283 net0513:F291 1918.19
R879 net0513:F267 net0513:F251 17288.8
R88 A:F163 A:F147 15098.7
R880 net0513:F251 net0513:F75 363.085
R881 net0513:F251 net0513:F71 1279.84
R882 net0513:F251 net0513:F67 4512.25
R883 net0513:F251 net0513:F63 15905.8
R884 net0513:F142 net0513:F182 705.36
R885 net0513:F142 net0513:F174 684.148
R886 net0513:F142 net0513:F166 646.526
R887 net0513:F142 net0513:F158 596.568
R888 net0513:F142 net0513:F150 746.745
R889 net0513:F142 net0513:F148 0.001
R89 A:F163 A:F3 130.382
R890 net0513:F150 net0513:F182 419.413
R891 net0513:F150 net0513:F174 406.801
R892 net0513:F150 net0513:F166 384.43
R893 net0513:F150 net0513:F158 354.725
R894 net0513:F150 net0513:F156 0.001
R895 net0513:F158 net0513:F182 298.747
R896 net0513:F158 net0513:F174 289.763
R897 net0513:F158 net0513:F166 273.829
R898 net0513:F158 net0513:F164 0.001
R899 net0513:F166 net0513:F182 226.756
R9 vdd vdd 0.001
R90 A:F167 A:F351 6774.68
R900 net0513:F166 net0513:F174 219.937
R901 net0513:F166 net0513:F172 0.001
R902 net0513:F174 net0513:F182 178.586
R903 net0513:F174 net0513:F180 0.001
R904 net0513:F31 net0513:F211 1280.37
R905 net0513:F31 net0513:F203 103.045
R906 net0513:F31 net0513:F195 1280.55
R907 net0513:F31 net0513:F187 10800.7
R908 net0513:F31 net0513:F47 15911.7
R909 net0513:F31 net0513:F43 4511.79
R91 A:F167 A:F347 2069.79
R910 net0513:F31 net0513:F39 1280.37
R911 net0513:F31 net0513:F35 357.956
R912 net0513:F31 net0513:F27 362.916
R913 net0513:F31 net0513:F23 1280.55
R914 net0513:F31 net0513:F19 3743.94
R915 net0513:F31 net0513:F15 10368.6
R916 net0513:F35 net0513:F211 363.222
R917 net0513:F35 net0513:F203 357.956
R918 net0513:F35 net0513:F195 4452.61
R919 net0513:F35 net0513:F187 19199.1
R92 A:F167 A:F343 446.147
R920 net0513:F35 net0513:F51 16007
R921 net0513:F35 net0513:F47 4513.92
R922 net0513:F35 net0513:F43 1279.93
R923 net0513:F35 net0513:F39 363.222
R924 net0513:F35 net0513:F27 1261.9
R925 net0513:F35 net0513:F23 4452.61
R926 net0513:F35 net0513:F19 15242.5
R927 net0513:F35 net0513:F15 18431.1
R928 net0513:F19 net0513:F203 4298.34
R929 net0513:F19 net0513:F195 345.745
R93 A:F167 A:F339 103.176
R930 net0513:F19 net0513:F187 265.731
R931 net0513:F19 net0513:F27 1218.8
R932 net0513:F19 net0513:F23 345.745
R933 net0513:F19 net0513:F15 255.101
R934 net0513:F39 net0513:F211 103.041
R935 net0513:F39 net0513:F203 1280.37
R936 net0513:F39 net0513:F195 13718.7
R937 net0513:F39 net0513:F59 24637
R938 net0513:F39 net0513:F55 13858.5
R939 net0513:F39 net0513:F51 4511.76
R94 A:F167 A:F335 379.921
R940 net0513:F39 net0513:F47 1279.88
R941 net0513:F39 net0513:F43 363.084
R942 net0513:F39 net0513:F27 3887.96
R943 net0513:F39 net0513:F23 13718.7
R944 net0513:F43 net0513:F211 363.084
R945 net0513:F43 net0513:F203 4511.79
R946 net0513:F43 net0513:F195 28061
R947 net0513:F43 net0513:F59 16007.6
R948 net0513:F43 net0513:F55 3931.48
R949 net0513:F43 net0513:F51 1279.93
R95 A:F167 A:F331 1873.03
R950 net0513:F43 net0513:F47 363.085
R951 net0513:F43 net0513:F27 15905.4
R952 net0513:F43 net0513:F23 28061
R953 net0513:F23 net0513:F211 15926.5
R954 net0513:F23 net0513:F203 1281.78
R955 net0513:F23 net0513:F195 103.155
R956 net0513:F23 net0513:F187 997.418
R957 net0513:F23 net0513:F27 363.623
R958 net0513:F23 net0513:F15 957.521
R959 net0513:F47 net0513:F211 1279.88
R96 A:F167 A:F327 4881.79
R960 net0513:F47 net0513:F203 15911.7
R961 net0513:F47 net0513:F67 24637.1
R962 net0513:F47 net0513:F63 13864
R963 net0513:F47 net0513:F59 4513.6
R964 net0513:F47 net0513:F55 1280.27
R965 net0513:F47 net0513:F51 363.22
R966 net0513:F27 net0513:F211 4513.67
R967 net0513:F27 net0513:F203 363.264
R968 net0513:F27 net0513:F195 363.623
R969 net0513:F27 net0513:F187 3516.04
R97 A:F167 A:F323 24183.1
R970 net0513:F27 net0513:F15 3375.4
R971 net0513:F51 net0513:F211 4511.76
R972 net0513:F51 net0513:F67 16008.1
R973 net0513:F51 net0513:F63 3933.16
R974 net0513:F51 net0513:F59 1280.49
R975 net0513:F51 net0513:F55 363.206
R976 net0513:F59 net0513:F211 24637
R977 net0513:F59 net0513:F75 16002.2
R978 net0513:F59 net0513:F71 3931.7
R979 net0513:F59 net0513:F67 1280.02
R98 A:F167 A:F179 7790.88
R980 net0513:F59 net0513:F63 363.236
R981 net0513:F59 net0513:F55 362.902
R982 net0513:F67 net0513:F75 1279.49
R983 net0513:F67 net0513:F71 363.087
R984 net0513:F67 net0513:F63 363.097
R985 net0513:F67 net0513:F55 4507.81
R986 net0513:F75 net0513:F71 363.084
R987 net0513:F75 net0513:F63 4510.22
R988 net0513:F75 net0513:F55 24605.5
R989 net0513:F55 net0513:F211 13858.5
R99 A:F167 A:F175 2380.26
R990 net0513:F55 net0513:F71 13846.2
R991 net0513:F55 net0513:F63 1279.2
R992 net0513:F63 net0513:F71 1279.89
R993 net0513:F187 net0513:F203 12400
R994 net0513:F187 net0513:F195 997.418
R995 net0513:F187 net0513:F15 77.2251
R996 net0513:F195 net0513:F211 15926.5
R997 net0513:F195 net0513:F203 1281.78
R998 net0513:F195 net0513:F15 957.521
R999 net0513:F203 net0513:F211 1280.37
.ENDS HS65_GS_BFX284


.SUBCKT HS65_GS_CB4I6X9 Z D C B A gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:12 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.212 PJ=7.32
MMM0 net072:F36 A:F37 gnd gnd NSVTGP AD=0.0561p AS=0.033p L=0.06u NRD=0.333333 NRS=0.333333 PD=0.67u PS=0.2u W=0.33u lpe=3 ngcon=1 po2act=0.288483 sca=3.10896 scb=0.00160583 scc=7.7901e-06
MMM1 net072:F34 B:F33 gnd gnd NSVTGP L=0.06u W=0.33u ad=0.033p as=0.033p lpe=3 ngcon=1 nrd=0.333333 nrs=0.333333 pd=0.2u po2act=0.51806 ps=0.2u sca=3.10862 scb=0.00160583 scc=7.7901e-06
MMM2 net050:F24 D:F25 gnd gnd NSVTGP AD=0.02332p AS=0.03113p L=0.06u NRD=0.25 NRS=0.643182 PD=0.204u PS=0.2222u W=0.22u lpe=3 ngcon=1 po2act=0.619858 sca=3.5329 scb=0.00216379 scc=1.15056e-05
MMM3 Z:F22 net050:F21 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.1365p as=0.11037p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=1.13u po2act=0.193633 ps=0.7878u sca=6.99153 scb=0.00671895 scc=0.000548722
MMM4 net050:F30 C:F29 net072:F28 gnd NSVTGP L=0.06u W=0.33u ad=0.03498p as=0.033p lpe=3 ngcon=1 nrd=0.333333 nrs=0.333333 pd=0.306u po2act=0.404915 ps=0.2u sca=3.1085 scb=0.00160583 scc=7.7901e-06
MMM5 net044:F44 D:F45 vdd vdd PSVTGP AD=0.066p AS=0.0713p L=0.06u NRD=0.490909 NRS=0.381818 PD=0.24u PS=0.333333u W=0.55u lpe=3 ngcon=1 po2act=0.619858 sca=2.376 scb=0.000974317 scc=4.28017e-06
MMM6 Z:F42 net050:F41 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.1925p as=0.1426p lpe=3 ngcon=1 nrd=0.25 nrs=0.295455 pd=1.45u po2act=0.217848 ps=0.666667u sca=5.22263 scb=0.00477169 scc=0.000389094
MMM7 net050:F54 B:F53 net048:F52 vdd PSVTGP L=0.06u W=0.55u ad=0.05775p as=0.04125p lpe=3 ngcon=1 nrd=0.327273 nrs=0.136364 pd=0.21u po2act=0.555177 ps=0.15u sca=2.37613 scb=0.000974317 scc=4.28017e-06
MMM8 net048:F58 A:F57 net044:F56 vdd PSVTGP L=0.06u W=0.55u ad=0.04125p as=0.0935p lpe=3 ngcon=1 nrd=0.136364 nrs=0.327273 pd=0.15u po2act=0.299007 ps=0.89u sca=2.37664 scb=0.000974317 scc=4.28017e-06
MMM9 net050:F48 C:F49 net044:F50 vdd PSVTGP AD=0.05775p AS=0.066p L=0.06u NRD=0.327273 NRS=0.327273 PD=0.21u PS=0.24u W=0.55u lpe=3 ngcon=1 po2act=0.700709 sca=2.37584 scb=0.000974317 scc=4.28017e-06
R1 net072:F28 net072:F36 76.0134
R10 A:F57 A:F37 322.366
R11 A:F57 A:F3 67.9433
R12 A:F3 A:F37 485.794
R13 net044:F50 net044:F56 76.0112
R14 net044:F50 net044:F44 0.001
R15 B B:F4 0.001
R16 B:F53 B:F4 171.834
R17 B:F53 B:F33 497.099
R18 B:F4 B:F33 186.898
R19 C C:F5 0.001
R2 net072:F28 net072:F34 0.001
R20 C:F49 C:F5 179.397
R21 C:F49 C:F29 489.603
R22 C:F5 C:F29 177.237
R23 D D:F6 0.001
R24 D:F45 D:F25 349.662
R25 D:F45 D:F6 432.753
R26 D:F6 D:F25 74.3862
R27 net050:F41 net050:F48 281.875
R28 net050:F41 net050:F24 279.869
R29 net050:F41 net050:F21 65.2582
R3 gnd gnd 0.001
R30 net050:F48 net050:F54 0.001
R31 net050:F48 net050:F24 107.826
R32 net050:F48 net050:F21 281.875
R33 net050:F21 net050:F24 279.869
R34 net050:F24 net050:F30 0.001
R35 Z Z:F7 0.001
R36 Z:F42 Z:F7 37.5
R37 Z:F7 Z:F22 38.4395
R38 vdd vdd 0.001
R39 vdd vdd 0.001
R4 gnd gnd 37.9799
R40 vdd vdd 0.001
R41 vdd vdd 0.001
R42 vdd vdd 0.001
R43 vdd vdd 0.001
R44 vdd vdd 37.6272
R45 vdd vdd 0.001
R46 vdd vdd 37.8033
R47 vdd vdd 0.001
R48 gnd gnd 0.001
R49 gnd gnd 0.001
R5 gnd gnd 37.6448
R50 gnd gnd 0.001
R51 gnd gnd 0.001
R52 gnd gnd 0.001
R53 gnd gnd 0.0256454
R54 gnd gnd 37.6257
R6 gnd gnd 0.001
R7 gnd gnd 0.001
R8 net048:F52 net048:F58 0.001
R9 A A:F3 0.001
.ENDS HS65_GS_CB4I6X9


.SUBCKT HS65_GS_CBI4I6X5 Z D C B A gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:12 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=2.92 PJ=6.92
MMM10 Z:F19 D:F20 gnd gnd NSVTGP AD=0.0484p AS=0.088p L=0.06u NRD=0.272727 NRS=0.136364 PD=0.256u PS=0.84u W=0.44u lpe=3 ngcon=1 po2act=0.333884 sca=5.80632 scb=0.00591115 scc=0.000194263
MMM11 Z:F25 C:F24 net033:F23 gnd NSVTGP L=0.06u W=0.66u ad=0.0726p as=0.0693p lpe=3 ngcon=1 nrd=0.272727 nrs=0.272727 pd=0.384u po2act=0.374961 ps=0.21u sca=4.53374 scb=0.00403577 scc=0.000129555
MMM12 net046:F47 B:F48 net93:F49 vdd PSVTGP AD=0.209p AS=0.121p L=0.06u NRD=0.272727 NRS=0.1 PD=1.48u PS=0.22u W=1.1u lpe=3 ngcon=1 po2act=0.320331 sca=5.22365 scb=0.00477169 scc=0.000389094
MMM13 net93:F43 A:F44 vdd vdd PSVTGP AD=0.121p AS=0.1155p L=0.06u NRD=0.1 NRS=0.272727 PD=0.22u PS=0.21u W=1.1u lpe=3 ngcon=1 po2act=0.574876 sca=5.22319 scb=0.00477169 scc=0.000389094
MMM14 net046:F41 C:F40 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.1155p as=0.1155p lpe=3 ngcon=1 nrd=0.272727 nrs=0.272727 pd=0.21u po2act=0.574876 ps=0.21u sca=5.22319 scb=0.00477169 scc=0.000389094
MMM2 Z:F37 D:F36 net046:F35 vdd PSVTGP L=0.06u W=1.1u ad=0.22p as=0.1155p lpe=3 ngcon=1 nrd=0.295455 nrs=0.272727 pd=1.5u po2act=0.333884 ps=0.21u sca=5.22363 scb=0.00477169 scc=0.000389094
MMM6 net033:F29 A:F28 gnd gnd NSVTGP L=0.06u W=0.66u ad=0.0693p as=0.0726p lpe=3 ngcon=1 nrd=0.272727 nrs=0.272727 pd=0.21u po2act=0.517881 ps=0.22u sca=4.53374 scb=0.00403577 scc=0.000129555
MMM9 net033:F31 B:F32 gnd gnd NSVTGP AD=0.1254p AS=0.0726p L=0.06u NRD=0.272727 NRS=0.318182 PD=1.04u PS=0.22u W=0.66u lpe=3 ngcon=1 po2act=0.312161 sca=4.53401 scb=0.00403577 scc=0.000129555
R1 net033:F23 net033:F31 75.6002
R10 B:F48 B:F32 107.313
R11 B:F48 B:F4 81.8576
R12 B:F4 B:F32 160.457
R13 A A:F3 0.001
R14 A:F44 A:F28 116.151
R15 A:F44 A:F3 84.6269
R16 A:F3 A:F28 159.937
R17 C C:F5 0.001
R18 C:F40 C:F24 116.077
R19 C:F40 C:F5 84.7396
R2 net033:F23 net033:F29 0.001
R20 C:F5 C:F24 160.15
R21 D D:F6 0.001
R22 D:F36 D:F20 105.987
R23 D:F36 D:F6 81.6055
R24 D:F6 D:F20 160.863
R25 Z Z:F7 0.001
R26 Z:F37 Z:F7 38.3857
R27 Z:F7 Z:F19 38.2317
R28 Z:F19 Z:F25 0.001
R29 vdd vdd 0.001
R3 gnd gnd 0.001
R30 vdd vdd 0.001
R31 vdd vdd 0.001
R32 vdd vdd 0.001
R33 vdd vdd 0.001
R34 vdd vdd 37.6252
R35 net93:F43 net93:F49 0.001
R36 vdd vdd 0.001
R37 vdd vdd 37.6461
R38 vdd vdd 0.001
R39 gnd gnd 0.001
R4 gnd gnd 37.688
R40 gnd gnd 0.001
R41 gnd gnd 0.001
R42 gnd gnd 0.001
R43 gnd gnd 0.0256454
R44 gnd gnd 37.6237
R5 gnd gnd 19.0727
R6 gnd gnd 0.001
R7 net046:F41 net046:F47 75.8729
R8 net046:F41 net046:F35 0.001
R9 B B:F4 0.001
.ENDS HS65_GS_CBI4I6X5


.SUBCKT HS65_GS_DFPQX4 Q D clk gnd gnd vdd vdd

*Modified
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:44 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=5.1312 PJ=10.24
MMM1 net47:F31R2 D gnd gnd NSVTGP AD=0.014p AS=0.0456667p L=0.06u NRD=0.35 NRS=0.4 PD=0.14u PS=0.530435u W=0.2u lpe=3 ngcon=1 po2act=0.296591 sca=1.69635 scb=0.000126319 scc=2.33728e-08
MMM12 R48 clk vdd vdd PSVTGP L=0.06u W=0.29u ad=0.058p as=0.0669495p lpe=3 ngcon=1 nrd=0.224138 nrs=15.3376 pd=0.69u po2act=0.28576 ps=0.636129u sca=14.0804 scb=0.0159942 scc=0.00146523
MMM13 R48 clk gnd gnd NSVTGP L=0.06u W=0.29u ad=0.05365p as=0.0662167p lpe=3 ngcon=1 nrd=0.206897 nrs=7.15869 pd=0.66u po2act=0.214753 ps=0.76913u sca=8.12641 scb=0.00955152 scc=0.000408996
MMM14 R32 R48 vdd vdd PSVTGP AD=0.0597p AS=0.0669495p L=0.06u NRD=0.344828 NRS=15.3376 PD=0.77u PS=0.636129u W=0.29u lpe=3 ngcon=1 po2act=0.275451 sca=14.0793 scb=0.0159942 scc=0.00146523
MMM15 R32 R48 gnd gnd NSVTGP AD=0.039p AS=0.0456667p L=0.06u NRD=0.3 NRS=8.2448 PD=0.59u PS=0.530435u W=0.2u lpe=3 ngcon=1 po2act=0.238627 sca=17.5984 scb=0.0199621 scc=0.00206349
MMM16 R27 R17 vdd vdd PSVTGP L=0.06u W=0.29u ad=0.0517p as=0.0623595p lpe=3 ngcon=1 nrd=0.206897 nrs=10.6859 pd=0.69u po2act=0.214968 ps=0.763158u sca=12.0121 scb=0.0141722 scc=0.00107611
MMM17 R27 R17 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.038p as=0.0500821p lpe=3 ngcon=1 nrd=0.3 nrs=10.1217 pd=0.58u po2act=0.326495 ps=0.564179u sca=17.5978 scb=0.0199621 scc=0.00206349
MMM18 net0109:F47R1 R27 gnd gnd NSVTGP AD=0.014p AS=0.0500821p L=0.06u NRD=0.35 NRS=2.20697 PD=0.14u PS=0.564179u W=0.2u lpe=3 ngcon=1 po2act=0.282173 sca=2.32991 scb=0.000604316 scc=6.73457e-07
MMM19 R17 R32 net0109:F47R1 gnd NSVTGP AD=0.035p AS=0.014p L=0.06u NRD=0.275 NRS=0.35 PD=0.55u PS=0.14u W=0.2u lpe=3 ngcon=1 po2act=0.24913 sca=2.33003 scb=0.000604316 scc=6.73457e-07
MMM20 R17 R48 net053:F103R12 vdd PSVTGP AD=0.037p AS=0.014p L=0.06u NRD=0.3 NRS=0.35 PD=0.57u PS=0.14u W=0.2u lpe=3 ngcon=1 po2act=0.247344 sca=1.54672 scb=0.000125995 scc=2.33727e-08
MMM21 net053:F103R12 R27 vdd vdd PSVTGP AD=0.014p AS=0.0430066p L=0.06u NRD=0.35 NRS=1.97518 PD=0.14u PS=0.526316u W=0.2u lpe=3 ngcon=1 po2act=0.23417 sca=1.54656 scb=0.000125995 scc=2.33727e-08
MMM22 R7 R27 vdd vdd PSVTGP AD=0.027p AS=0.0580589p L=0.06u NRD=0.203704 NRS=10.8032 PD=0.2u PS=0.710526u W=0.27u lpe=3 ngcon=1 po2act=0.373692 sca=6.20515 scb=0.00679075 scc=0.000173611
MMM23 R7 R27 gnd gnd NSVTGP AD=0.029025p AS=0.0676108p L=0.06u NRD=0.240741 NRS=9.38888 PD=0.215u PS=0.761642u W=0.27u lpe=3 ngcon=1 po2act=0.454622 sca=14.7788 scb=0.0167784 scc=0.00156883
MMM24 R7 R48 R62 vdd PSVTGP L=0.06u W=0.27u ad=0.027p as=0.0347266p lpe=3 ngcon=1 nrd=0.203704 nrs=0.333333 pd=0.2u po2act=0.371244 ps=0.373404u sca=6.20538 scb=0.00679075 scc=0.000173611
MMM25 R7 R32 R62 gnd NSVTGP L=0.06u W=0.27u ad=0.029025p as=0.0322071p lpe=3 ngcon=1 nrd=0.222222 nrs=0.259259 pd=0.215u po2act=0.363522 ps=0.372857u sca=14.779 scb=0.0167784 scc=0.00156883
MMM26 net069:F115R4 R39 vdd vdd PSVTGP L=0.06u W=0.2u ad=0.017p as=0.0364737p lpe=3 ngcon=1 nrd=0.425 nrs=8.68125 pd=0.17u po2act=0.630845 ps=0.349474u sca=6.20704 scb=0.00684993 scc=0.000149357
MMM27 R62 R32 net069:F115R4 vdd PSVTGP L=0.06u W=0.2u ad=0.0257234p as=0.017p lpe=3 ngcon=1 nrd=0.375 nrs=0.425 pd=0.276596u po2act=0.571307 ps=0.17u sca=8.55791 scb=0.0105547 scc=0.000414651
MMM28 R39 R62 vdd vdd PSVTGP L=0.06u W=0.2u ad=0.082425p as=0.0364737p lpe=3 ngcon=1 nrd=1.74938 nrs=0.3 pd=1.13u po2act=0.211059 ps=0.349474u sca=1.10977 scb=1.22045e-05 scc=1.68552e-10
MMM29 R62 R48 net0133:F63R3 gnd NSVTGP L=0.06u W=0.15u ad=0.0178929p as=0.0105p lpe=3 ngcon=1 nrd=0.466667 nrs=0.466667 pd=0.207143u po2act=0.820147 ps=0.14u sca=12.5289 scb=0.0158913 scc=0.00101939
MMM30 net0133:F63R3 R39 gnd gnd NSVTGP L=0.06u W=0.15u ad=0.0105p as=0.0273851p lpe=3 ngcon=1 nrd=0.466667 nrs=9.42667 pd=0.14u po2act=0.687885 ps=0.316216u sca=20.4056 scb=0.0226819 scc=0.00260982
MMM31 R39 R62 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0755p as=0.0365135p lpe=3 ngcon=1 nrd=1.7 nrs=0.35 pd=1.06u po2act=0.214984 ps=0.421622u sca=1.88439 scb=0.000214041 scc=7.20983e-08
MMM32 Q R62 vdd vdd PSVTGP AD=0.09075p AS=0.100303p L=0.06u NRD=0.3 NRS=6.18099 PD=0.88u PS=0.961053u W=0.55u lpe=3 ngcon=1 po2act=0.200385 sca=3.81818 scb=0.00308337 scc=5.58864e-05
MMM33 Q R62 gnd gnd NSVTGP AD=0.06435p AS=0.0712014p L=0.06u NRD=0.282051 NRS=6.64323 PD=0.72u PS=0.822162u W=0.39u lpe=3 ngcon=1 po2act=0.192123 sca=11.6369 scb=0.0127786 scc=0.00109616
MMM4 R17 R48 net47:F31R2 gnd NSVTGP AD=0.0862p AS=0.014p L=0.06u NRD=1.78633 NRS=0.35 PD=1.16u PS=0.14u W=0.2u lpe=3 ngcon=1 po2act=0.302652 sca=1.69604 scb=0.000126319 scc=2.33728e-08
MMM5 R17 R32 net22:F81R36 vdd PSVTGP AD=0.0612p AS=0.0558p L=0.06u NRD=0.323529 NRS=0.323529 PD=0.7u PS=0.7u W=0.34u lpe=3 ngcon=1 po2act=0.17 sca=1.72715 scb=0.000243274 scc=1.32953e-07
MMM6 net22:F81R36 D vdd vdd PSVTGP L=0.06u W=0.35u ad=0.05775p as=0.0808011p lpe=3 ngcon=1 nrd=0.314286 nrs=0.885714 pd=0.68u po2act=0.211816 ps=0.767742u sca=1.36111 scb=6.68153e-05 scc=8.8344e-09


.ENDS HS65_GS_DFPQX4


.SUBCKT HS65_GS_DFPQX9 Q D CP gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:44 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=5.1312 PJ=10.24
MMM1 net47:F31 D:F32 gnd gnd NSVTGP AD=0.014p AS=0.0456667p L=0.06u NRD=0.35 NRS=0.4 PD=0.14u PS=0.530435u W=0.2u lpe=3 ngcon=1 po2act=0.296591 sca=1.69635 scb=0.000126319 scc=2.33728e-08
MMM12 CPN:F85 CP:F84 vdd vdd PSVTGP L=0.06u W=0.29u ad=0.058p as=0.0669495p lpe=3 ngcon=1 nrd=0.224138 nrs=15.3376 pd=0.69u po2act=0.28576 ps=0.636129u sca=14.0804 scb=0.0159942 scc=0.00146523
MMM13 CPN:F29 CP:F28 gnd gnd NSVTGP L=0.06u W=0.29u ad=0.05365p as=0.0662167p lpe=3 ngcon=1 nrd=0.206897 nrs=7.15869 pd=0.66u po2act=0.214904 ps=0.76913u sca=8.12641 scb=0.00955152 scc=0.000408996
MMM14 CPI:F87 CPN:F88 vdd vdd PSVTGP AD=0.0597p AS=0.0669495p L=0.06u NRD=0.344828 NRS=15.3376 PD=0.77u PS=0.636129u W=0.29u lpe=3 ngcon=1 po2act=0.275451 sca=14.0793 scb=0.0159942 scc=0.00146523
MMM15 CPI:F35 CPN:F36 gnd gnd NSVTGP AD=0.04p AS=0.0456667p L=0.06u NRD=0.35 NRS=8.2448 PD=0.6u PS=0.530435u W=0.2u lpe=3 ngcon=1 po2act=0.242334 sca=17.5984 scb=0.0199621 scc=0.00206349
MMM16 net0113:F97 net35:F96 vdd vdd PSVTGP L=0.06u W=0.29u ad=0.0517p as=0.0623595p lpe=3 ngcon=1 nrd=0.189655 nrs=10.6859 pd=0.69u po2act=0.214968 ps=0.763158u sca=12.0121 scb=0.0141722 scc=0.00107611
MMM17 net0113:F45 net35:F44 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.04p as=0.0500821p lpe=3 ngcon=1 nrd=0.35 nrs=10.1217 pd=0.6u po2act=0.34039 ps=0.564179u sca=17.5978 scb=0.0199621 scc=0.00206349
MMM18 net0109:F47 net0113:F48 gnd gnd NSVTGP AD=0.014p AS=0.0500821p L=0.06u NRD=0.35 NRS=2.20697 PD=0.14u PS=0.564179u W=0.2u lpe=3 ngcon=1 po2act=0.283577 sca=2.32992 scb=0.000604316 scc=6.73457e-07
MMM19 net35:F55 CPI:F56 net0109:F57 gnd NSVTGP AD=0.036p AS=0.014p L=0.06u NRD=0.275 NRS=0.35 PD=0.56u PS=0.14u W=0.2u lpe=3 ngcon=1 po2act=0.254156 sca=2.33005 scb=0.000604316 scc=6.73457e-07
MMM20 net35:F107 CPN:F108 net053:F109 vdd PSVTGP AD=0.038p AS=0.014p L=0.06u NRD=0.275 NRS=0.35 PD=0.58u PS=0.14u W=0.2u lpe=3 ngcon=1 po2act=0.251773 sca=1.54672 scb=0.000125995 scc=2.33727e-08
MMM21 net053:F103 net0113:F104 vdd vdd PSVTGP AD=0.014p AS=0.0430066p L=0.06u NRD=0.35 NRS=1.97518 PD=0.14u PS=0.526316u W=0.2u lpe=3 ngcon=1 po2act=0.235087 sca=1.54656 scb=0.000125995 scc=2.33727e-08
MMM22 net0145:F99 net0113:F100 vdd vdd PSVTGP AD=0.027p AS=0.0580589p L=0.06u NRD=0.203704 NRS=10.8032 PD=0.2u PS=0.710526u W=0.27u lpe=3 ngcon=1 po2act=0.373692 sca=6.20515 scb=0.00679075 scc=0.000173611
MMM23 net0145:F51 net0113:F52 gnd gnd NSVTGP AD=0.027p AS=0.0676108p L=0.06u NRD=0.203704 NRS=9.38888 PD=0.2u PS=0.761642u W=0.27u lpe=3 ngcon=1 po2act=0.452589 sca=14.7788 scb=0.0167784 scc=0.00156883
MMM24 net0145:F113 CPN:F112 net0148:F111 vdd PSVTGP L=0.06u W=0.27u ad=0.027p as=0.0347266p lpe=3 ngcon=1 nrd=0.203704 nrs=0.333333 pd=0.2u po2act=0.371244 ps=0.373404u sca=6.20538 scb=0.00679075 scc=0.000173611
MMM25 net0145:F61 CPI:F60 net0148:F59 gnd NSVTGP L=0.06u W=0.27u ad=0.027p as=0.0322071p lpe=3 ngcon=1 nrd=0.203704 nrs=0.203704 pd=0.2u po2act=0.361874 ps=0.372857u sca=14.779 scb=0.0167784 scc=0.00156883
MMM26 net069:F121 net097:F120 vdd vdd PSVTGP L=0.06u W=0.2u ad=0.014p as=0.02784p lpe=3 ngcon=1 nrd=0.35 nrs=0.696 pd=0.14u po2act=0.642131 ps=0.202667u sca=6.20693 scb=0.00684993 scc=0.000149357
MMM27 net0148:F117 CPI:F116 net069:F115 vdd PSVTGP L=0.06u W=0.2u ad=0.0257234p as=0.014p lpe=3 ngcon=1 nrd=0.375 nrs=0.35 pd=0.276596u po2act=0.571307 ps=0.14u sca=8.55791 scb=0.0105547 scc=0.000414651
MMM28 net097:F125 net0148:F124 vdd vdd PSVTGP L=0.06u W=0.2u ad=0.0856p as=0.02784p lpe=3 ngcon=1 nrd=1.7625 nrs=0.425 pd=1.15u po2act=0.318881 ps=0.202667u sca=1.10984 scb=1.22045e-05 scc=1.68552e-10
MMM29 net0148:F65 CPN:F64 net0133:F63 gnd NSVTGP L=0.06u W=0.15u ad=0.0178929p as=0.0105p lpe=3 ngcon=1 nrd=0.566667 nrs=0.466667 pd=0.207143u po2act=0.818177 ps=0.14u sca=12.5289 scb=0.0158913 scc=0.00101939
MMM30 net0133:F69 net097:F68 gnd gnd NSVTGP L=0.06u W=0.15u ad=0.0105p as=0.017708p lpe=3 ngcon=1 nrd=0.466667 nrs=0.787021 pd=0.14u po2act=0.686938 ps=0.142035u sca=20.4056 scb=0.0226819 scc=0.00260982
MMM31 net097:F73 net0148:F72 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.07225p as=0.0236106p lpe=3 ngcon=1 nrd=1.62667 nrs=0.275 pd=1.03u po2act=0.272 ps=0.189381u sca=1.88439 scb=0.000214041 scc=7.20983e-08
MMM32 Q:F127 net0148:F128 vdd vdd PSVTGP AD=0.1815p AS=0.15312p L=0.06u NRD=0.25 NRS=0.340909 PD=1.43u PS=1.11467u W=1.1u lpe=3 ngcon=1 po2act=0.181115 sca=5.21719 scb=0.00477169 scc=0.000389094
MMM33 Q:F75 net0148:F76 gnd gnd NSVTGP AD=0.1287p AS=0.0920814p L=0.06u NRD=0.282051 NRS=0.282051 PD=1.11u PS=0.738584u W=0.78u lpe=3 ngcon=1 po2act=0.182107 sca=6.98771 scb=0.00671895 scc=0.000548722
MMM4 net35:F39 CPN:F40 net47:F41 gnd NSVTGP AD=0.0862p AS=0.014p L=0.06u NRD=1.78633 NRS=0.35 PD=1.16u PS=0.14u W=0.2u lpe=3 ngcon=1 po2act=0.302652 sca=1.69604 scb=0.000126319 scc=2.33728e-08
MMM5 net35:F91 CPI:F92 net22:F93 vdd PSVTGP AD=0.0612p AS=0.0558p L=0.06u NRD=0.323529 NRS=0.323529 PD=0.7u PS=0.7u W=0.34u lpe=3 ngcon=1 po2act=0.17 sca=1.72715 scb=0.000243274 scc=1.32953e-07
MMM6 net22:F81 D:F80 vdd vdd PSVTGP L=0.06u W=0.35u ad=0.05775p as=0.0808011p lpe=3 ngcon=1 nrd=0.314286 nrs=0.885714 pd=0.68u po2act=0.211816 ps=0.767742u sca=1.36111 scb=6.68153e-05 scc=8.8344e-09
R1 net0109:F47 net0109:F57 0.001
R10 CP:F84 CP:F28 108.835
R100 gnd gnd 0.001
R101 gnd gnd 0.001
R102 gnd gnd 0.001
R103 gnd gnd 0.001
R104 gnd gnd 0.001
R105 gnd gnd 0.001
R106 gnd gnd 0.001
R107 gnd gnd 0.001
R108 gnd gnd 0.001
R109 gnd gnd 0.001
R11 CP:F3 CP:F28 149.773
R110 gnd gnd 3412.5
R111 gnd gnd 2680.16
R112 gnd gnd 3368.01
R113 gnd gnd 2.17112
R114 gnd gnd 38.7753
R115 gnd gnd 38.7053
R116 gnd gnd 38.2697
R117 gnd gnd 6332.96
R118 gnd gnd 0.001
R119 gnd gnd 0.001
R12 net053:F103 net053:F109 0.001
R120 gnd gnd 0.001
R121 gnd gnd 0.001
R122 gnd gnd 0.001
R123 gnd gnd 0.001
R13 net35:F91 net35:F107 89.345
R14 net35:F91 net35:F96 252.277
R15 net35:F107 net35:F96 255.955
R16 net35:F96 net35:F44 79
R17 net35:F44 net35:F39 191.322
R18 net35:F44 net35:F55 194.76
R19 net35:F39 net35:F55 94.7159
R2 net0133:F63 net0133:F69 0.001
R20 net0113:F104 net0113:F100 58.75
R21 net0113:F100 net0113:F97 359.131
R22 net0113:F100 net0113:F52 120.87
R23 net0113:F100 net0113:F45 362.072
R24 net0113:F97 net0113:F52 277.47
R25 net0113:F97 net0113:F45 99.6942
R26 net0113:F52 net0113:F45 279.742
R27 net0113:F52 net0113:F48 47.5
R28 CPI:F92 CPI:F116 308.263
R29 CPI:F92 CPI:F87 185.825
R3 net47:F31 net47:F41 0.001
R30 CPI:F92 CPI:F35 187.576
R31 CPI:F116 CPI:F87 206.802
R32 CPI:F116 CPI:F60 159.5
R33 CPI:F116 CPI:F35 208.751
R34 CPI:F87 CPI:F35 125.838
R35 CPI:F60 CPI:F56 36.25
R36 net22:F81 net22:F93 75.8084
R37 net097:F125 net097:F120 99.0947
R38 net097:F68 net097:F120 114.081
R39 net097:F68 net097:F73 161.52
R4 net069:F115 net069:F121 0.001
R40 net097:F120 net097:F73 245.145
R41 net0148:F128 net0148:F124 132.5
R42 net0148:F128 net0148:F111 284.058
R43 net0148:F128 net0148:F76 70.1696
R44 net0148:F128 net0148:F59 290.255
R45 net0148:F111 net0148:F117 0.001
R46 net0148:F111 net0148:F76 284.058
R47 net0148:F111 net0148:F59 103.018
R48 net0148:F76 net0148:F72 120
R49 net0148:F76 net0148:F59 290.255
R5 net0145:F99 net0145:F113 0.001
R50 net0148:F59 net0148:F65 0.001
R51 CPN:F108 CPN:F112 48.125
R52 CPN:F108 CPN:F88 567.75
R53 CPN:F88 CPN:F85 277.006
R54 CPN:F88 CPN:F36 61.8276
R55 CPN:F88 CPN:F29 278.887
R56 CPN:F85 CPN:F36 277.006
R57 CPN:F85 CPN:F29 106.356
R58 CPN:F36 CPN:F40 148.75
R59 CPN:F36 CPN:F29 278.887
R6 net0145:F99 net0145:F51 75.9438
R60 CPN:F64 CPN:F40 516.25
R61 D D:F4 0.001
R62 D:F80 D:F32 3615.3
R63 D:F80 D:F4 310.38
R64 D:F4 D:F32 540.463
R65 Q Q:F5 0.001
R66 Q:F5 Q:F127 37.6364
R67 Q:F5 Q:F75 38.6369
R68 vdd vdd 0.001
R69 vdd vdd 38.4288
R7 net0145:F51 net0145:F61 0.001
R70 vdd vdd 38.1366
R71 vdd vdd 37.5667
R72 vdd vdd 0.001
R73 vdd vdd 0.001
R74 vdd vdd 0.001
R75 vdd vdd 0.001
R76 vdd vdd 4510.34
R77 vdd vdd 0.001
R78 vdd vdd 0.001
R79 vdd vdd 0.001
R8 CP CP:F3 0.001
R80 vdd vdd 0.001
R81 vdd vdd 0.001
R82 vdd vdd 0.001
R83 vdd vdd 0.001
R84 vdd vdd 0.001
R85 vdd vdd 0.001
R86 vdd vdd 0.001
R87 vdd vdd 0.001
R88 vdd vdd 0.001
R89 vdd vdd 0.001
R9 CP:F84 CP:F3 86.377
R90 vdd vdd 0.001
R91 vdd vdd 0.001
R92 vdd vdd 0.001
R93 vdd vdd 37.6257
R94 gnd gnd 0.001
R95 gnd gnd 0.0256454
R96 gnd gnd 37.6237
R97 gnd gnd 0.001
R98 gnd gnd 0.001
R99 gnd gnd 0.001
.ENDS HS65_GS_DFPQX9


.SUBCKT HS65_GS_IVX9 Z A gnd gnd vdd vdd
*Modified

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:17 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=1.752 PJ=5.32
MMM64 Z:F13 A:F14 gnd gnd NSVTGP AD=0.1599p AS=0.1599p L=0.06u NRD=0.358974 NRS=0.358974 PD=1.19u PS=1.19u W=0.78u lpe=3 ngcon=1 po2act=0.205 sca=6.99573 scb=0.00671895 scc=0.000548722
MMM65 Z:F17 A:F18 vdd vdd PSVTGP AD=0.2255p AS=0.2255p L=0.06u NRD=0.159091 NRS=0.318182 PD=1.51u PS=1.51u W=1.1u lpe=3 ngcon=1 po2act=0.205 sca=5.22897 scb=0.00477169 scc=0.000389094
R1 gnd gnd 0.001
R10 vdd vdd 0.001
R11 vdd vdd 0.001
R12 vdd vdd 37.6252
R13 vdd vdd 0.001
R14 vdd vdd 37.5134
R15 gnd gnd 0.001
R16 gnd gnd 0.0256454
R17 gnd gnd 37.6237
R2 gnd gnd 37.5194
R3 Z Z:F4 0.001
R4 Z:F17 Z:F4 19.2183
R5 Z:F4 Z:F13 37.6912
R6 A A:F3 0.001
R7 A:F18 A:F14 71.6302
R8 A:F18 A:F3 101.631
R9 A:F3 A:F14 101.631
.ENDS HS65_GS_IVX9


.SUBCKT HS65_GS_MUX21X4 D0 D1 S0 Z gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:49 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.212 PJ=7.32
MMMN10 Z:F21 net16:F20 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.06435p as=0.0728441p lpe=3 ngcon=1 nrd=0.282051 nrs=4.78853 pd=0.72u po2act=0.198129 ps=0.932034u sca=11.6407 scb=0.0127786 scc=0.00109616
MMMN12 net8:F23 D0:F24 gnd gnd NSVTGP AD=0.02p AS=0.0373559p L=0.06u NRD=0.275 NRS=6.0175 PD=0.2u PS=0.477966u W=0.2u lpe=3 ngcon=1 po2act=0.512777 sca=9.16276 scb=0.0113099 scc=0.00048992
MMMN13 net5:F41 D1:F40 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0205p as=0.0707p lpe=3 ngcon=1 nrd=0.275 nrs=3.14444 pd=0.205u po2act=0.230588 ps=1.015u sca=17.6154 scb=0.0199621 scc=0.00206349
MMMN14 net8:F29 net20:F28 net16:F27 gnd NSVTGP L=0.06u W=0.2u ad=0.02p as=0.0296p lpe=3 ngcon=1 nrd=0.275 nrs=0.3 pd=0.2u po2act=0.441875 ps=0.35u sca=9.16263 scb=0.0113099 scc=0.00048992
MMMN15 net5:F35 S0:F36 net16:F37 gnd NSVTGP AD=0.0205p AS=0.0296p L=0.06u NRD=0.3 NRS=0.164543 PD=0.205u PS=0.35u W=0.2u lpe=3 ngcon=1 po2act=0.326806 sca=17.615 scb=0.0199621 scc=0.00206349
MMMN16 net20:F33 S0:F32 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.066p as=0.0707p lpe=3 ngcon=1 nrd=1.38333 nrs=0.35 pd=0.94u po2act=0.276585 ps=1.015u sca=1.95003 scb=0.000254845 scc=1.04822e-07
MMMP12 Z:F45 net16:F44 vdd vdd PSVTGP L=0.06u W=0.55u ad=0.09075p as=0.120975p lpe=3 ngcon=1 nrd=0.3 nrs=14.864 pd=0.88u po2act=0.19041 ps=1.085u sca=9.01084 scb=0.00942268 scc=0.00077814
MMMP14 net8:F47 D0:F48 vdd vdd PSVTGP AD=0.0475p AS=0.0615873p L=0.06u NRD=0.196429 NRS=15.7759 PD=0.545u PS=0.552364u W=0.28u lpe=3 ngcon=1 po2act=0.247917 sca=14.3941 scb=0.0163798 scc=0.00151539
MMMP15 net5:F65 D1:F64 vdd vdd PSVTGP L=0.06u W=0.28u ad=0.0307p as=0.11785p lpe=3 ngcon=1 nrd=0.196429 nrs=4.40741 pd=0.29u po2act=0.181404 ps=2.13u sca=6.58221 scb=0.00738115 scc=0.00021642
MMMP16 net8:F53 S0:F52 net16:F51 vdd PSVTGP L=0.06u W=0.28u ad=0.0475p as=0.03745p lpe=3 ngcon=1 nrd=5.83571 nrs=0.196429 pd=0.545u po2act=0.199902 ps=0.35u sca=2.97422 scb=0.00155102 scc=6.37382e-06
MMMP17 net5:F59 net20:F60 net16:F61 vdd PSVTGP AD=0.0307p AS=0.03745p L=0.06u NRD=0.196429 NRS=0.0623178 PD=0.29u PS=0.35u W=0.28u lpe=3 ngcon=1 po2act=0.234188 sca=4.37428 scb=0.00374731 scc=4.55614e-05
MMMP18 net20:F55 S0:F56 vdd vdd PSVTGP AD=0.0891p AS=0.0593877p L=0.06u NRD=1.05093 NRS=0.259259 PD=1.01u PS=0.532636u W=0.27u lpe=3 ngcon=1 po2act=0.317518 sca=1.15705 scb=1.85943e-05 scc=4.82094e-10
R1 gnd gnd 0.001
R10 D1 D1:F4 0.001
R11 D1:F64 D1:F4 112.532
R12 D1:F64 D1:F40 129.813
R13 D1:F4 D1:F40 122.465
R14 net5:F59 net5:F65 0.001
R15 net5:F59 net5:F41 76.8221
R16 net5:F41 net5:F35 0.001
R17 Z Z:F6 0.001
R18 Z:F45 Z:F6 37.7087
R19 Z:F6 Z:F21 37.8853
R2 gnd gnd 0.001
R20 net16:F44 net16:F51 148.659
R21 net16:F44 net16:F37 155.253
R22 net16:F44 net16:F20 70
R23 net16:F51 net16:F61 0.001
R24 net16:F51 net16:F37 103.003
R25 net16:F37 net16:F27 0.001
R26 net20:F55 net20:F60 249.248
R27 net20:F55 net20:F33 121.28
R28 net20:F55 net20:F28 199.895
R29 net20:F60 net20:F33 277.97
R3 gnd gnd 37.5761
R30 net20:F60 net20:F28 458.154
R31 net20:F28 net20:F33 178.646
R32 net8:F53 net8:F47 0.001
R33 net8:F53 net8:F29 76.1636
R34 net8:F29 net8:F23 0.001
R35 S0 S0:F5 0.001
R36 S0:F56 S0:F5 143.959
R37 S0:F56 S0:F52 46.4537
R38 S0:F5 S0:F52 143.959
R39 S0:F52 S0:F36 216.083
R4 gnd gnd 0.001
R40 S0:F36 S0:F32 90
R41 vdd vdd 0.001
R42 vdd vdd 0.001
R43 vdd vdd 0.001
R44 vdd vdd 0.001
R45 vdd vdd 0.001
R46 vdd vdd 0.001
R47 vdd vdd 0.001
R48 vdd vdd 37.6272
R49 vdd vdd 0.001
R5 gnd gnd 19.0799
R50 vdd vdd 37.8278
R51 vdd vdd 18.9624
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 gnd gnd 0.001
R55 gnd gnd 0.001
R56 gnd gnd 0.001
R57 gnd gnd 0.001
R58 gnd gnd 0.001
R59 gnd gnd 0.001
R6 D0 D0:F3 0.001
R60 gnd gnd 0.0256454
R61 gnd gnd 37.6257
R7 D0:F48 D0:F3 85.3073
R8 D0:F48 D0:F24 112.618
R9 D0:F3 D0:F24 156.023
.ENDS HS65_GS_MUX21X4


.SUBCKT HS65_GS_MUX21X44 D0 D1 S0 Z gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070516.0 at 17:52 5 Jun 2007
Xld_D0 gnd vdd DNWPS AREA=9.052 PJ=15.32
MMMN10 Z:F75 net16:F76 gnd gnd NSVTGP AD=0.078p AS=0.0812453p L=0.06u NRD=0.141026 NRS=0.282051 PD=0.2u PS=0.335912u W=0.78u lpe=3 ngcon=1 po2act=0.668091 sca=6.9826 scb=0.00671895 scc=0.000548722
MMMN10@2 Z:F81 net16:F80 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.282051 pd=0.2u po2act=1.03181 ps=0.2u sca=6.98355 scb=0.00671895 scc=0.000548722
MMMN10@3 Z:F83 net16:F84 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.141026 NRS=0.282051 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=0.97459 sca=6.9846 scb=0.00671895 scc=0.000548722
MMMN10@4 Z:F89 net16:F88 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.141026 nrs=0.282051 pd=0.2u po2act=0.72212 ps=0.2u sca=6.98575 scb=0.00671895 scc=0.000548722
MMMN10@5 Z:F91 net16:F92 gnd gnd NSVTGP AD=0.1404p AS=0.078p L=0.06u NRD=0.153846 NRS=0.282051 PD=1.14u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=0.334659 sca=6.98703 scb=0.00671895 scc=0.000548722
MMMN12 net8:F21 D0:F20 gnd gnd NSVTGP L=0.06u W=0.59u ad=0.1062p as=0.06195p lpe=3 ngcon=1 nrd=0.305085 nrs=0.305085 pd=0.95u po2act=0.310603 ps=0.21u sca=8.6356 scb=0.00881748 scc=0.000725408
MMMN12@2 net8:F23 D0:F24 gnd gnd NSVTGP AD=0.06195p AS=0.06195p L=0.06u NRD=0.305085 NRS=0.305085 PD=0.21u PS=0.21u W=0.59u lpe=3 ngcon=1 po2act=0.589714 sca=8.63427 scb=0.00881748 scc=0.000725408
MMMN12@3 net8:F29 D0:F28 gnd gnd NSVTGP L=0.06u W=0.59u ad=0.06195p as=0.06195p lpe=3 ngcon=1 nrd=0.305085 nrs=0.305085 pd=0.21u po2act=0.637989 ps=0.21u sca=8.63308 scb=0.00881748 scc=0.000725408
MMMN13 net5:F65 D1:F64 gnd gnd NSVTGP L=0.06u W=0.59u ad=0.059p as=0.059p lpe=3 ngcon=1 nrd=0.279661 nrs=0.279661 pd=0.2u po2act=1.86096 ps=0.2u sca=8.6288 scb=0.00881748 scc=0.000725408
MMMN13@2 net5:F67 D1:F68 gnd gnd NSVTGP AD=0.059p AS=0.059p L=0.06u NRD=0.279661 NRS=0.279661 PD=0.2u PS=0.2u W=0.59u lpe=3 ngcon=1 po2act=1.86096 sca=8.62952 scb=0.00881748 scc=0.000725408
MMMN13@3 net5:F73 D1:F72 gnd gnd NSVTGP L=0.06u W=0.59u ad=0.059p as=0.0614547p lpe=3 ngcon=1 nrd=0.279661 nrs=0.279661 pd=0.2u po2act=1.78866 ps=0.254088u sca=8.63031 scb=0.00881748 scc=0.000725408
MMMN14 net8:F41 net20:F40 net16:F39 gnd NSVTGP L=0.06u W=0.59u ad=0.1062p as=0.059p lpe=3 ngcon=1 nrd=0.305085 nrs=0.279661 pd=0.95u po2act=0.342674 ps=0.2u sca=8.62921 scb=0.00881748 scc=0.000725408
MMMN14@2 net8:F43 net20:F44 net16:F45 gnd NSVTGP AD=0.059p AS=0.059p L=0.06u NRD=0.279661 NRS=0.279661 PD=0.2u PS=0.2u W=0.59u lpe=3 ngcon=1 po2act=0.776471 sca=8.62851 scb=0.00881748 scc=0.000725408
MMMN14@3 net8:F49 net20:F48 net16:F47 gnd NSVTGP L=0.06u W=0.59u ad=0.059p as=0.059p lpe=3 ngcon=1 nrd=0.279661 nrs=0.279661 pd=0.2u po2act=1.13797 ps=0.2u sca=8.62787 scb=0.00881748 scc=0.000725408
MMMN15 net5:F51 S0:F52 net16:F53 gnd NSVTGP AD=0.059p AS=0.059p L=0.06u NRD=0.279661 NRS=0.279661 PD=0.2u PS=0.2u W=0.59u lpe=3 ngcon=1 po2act=1.42717 sca=8.6276 scb=0.00881748 scc=0.000725408
MMMN15@2 net5:F57 S0:F56 net16:F55 gnd NSVTGP L=0.06u W=0.59u ad=0.059p as=0.059p lpe=3 ngcon=1 nrd=0.279661 nrs=0.279661 pd=0.2u po2act=1.64406 ps=0.2u sca=8.62761 scb=0.00881748 scc=0.000725408
MMMN15@3 net5:F59 S0:F60 net16:F61 gnd NSVTGP AD=0.059p AS=0.059p L=0.06u NRD=0.279661 NRS=0.279661 PD=0.2u PS=0.2u W=0.59u lpe=3 ngcon=1 po2act=1.78866 sca=8.62813 scb=0.00881748 scc=0.000725408
MMMN16 net20:F31 S0:F32 gnd gnd NSVTGP AD=0.0838456p AS=0.06195p L=0.06u NRD=0.305085 NRS=0.305085 PD=0.511333u PS=0.21u W=0.59u lpe=3 ngcon=1 po2act=0.423825 sca=8.63201 scb=0.00881748 scc=0.000725408
MMMN16@2 net20:F37 S0:F36 gnd gnd NSVTGP L=0.06u W=0.31u ad=0.0440544p as=0.0558p lpe=3 ngcon=1 nrd=0.458423 nrs=0.193548 pd=0.268667u po2act=0.316216 ps=0.67u sca=3.36713 scb=0.00198702 scc=1.18733e-05
MMMP12 Z:F151 net16:F152 vdd vdd PSVTGP AD=0.11p AS=0.114813p L=0.06u NRD=0.125 NRS=0.25 PD=0.2u PS=0.389583u W=1.1u lpe=3 ngcon=1 po2act=0.650718 sca=5.20721 scb=0.00477169 scc=0.000389094
MMMP12@2 Z:F157 net16:F156 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.25 pd=0.2u po2act=1.01911 ps=0.2u sca=5.20861 scb=0.00477169 scc=0.000389094
MMMP12@3 Z:F159 net16:F160 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=0.968338 sca=5.21018 scb=0.00477169 scc=0.000389094
MMMP12@4 Z:F165 net16:F164 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.25 pd=0.2u po2act=0.719854 ps=0.2u sca=5.21194 scb=0.00477169 scc=0.000389094
MMMP12@5 Z:F167 net16:F168 vdd vdd PSVTGP AD=0.198p AS=0.11p L=0.06u NRD=0.136364 NRS=0.25 PD=1.46u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=0.334308 sca=5.21392 scb=0.00477169 scc=0.000389094
MMMP14 net8:F97 D0:F96 vdd vdd PSVTGP L=0.06u W=0.82u ad=0.1476p as=0.0861p lpe=3 ngcon=1 nrd=0.292683 nrs=0.292683 pd=1.18u po2act=0.307147 ps=0.21u sca=2.082 scb=0.000807962 scc=4.50361e-06
MMMP14@2 net8:F99 D0:F100 vdd vdd PSVTGP AD=0.0861p AS=0.0861p L=0.06u NRD=0.292683 NRS=0.292683 PD=0.21u PS=0.21u W=0.82u lpe=3 ngcon=1 po2act=0.557735 sca=2.07994 scb=0.000807962 scc=4.50361e-06
MMMP14@3 net8:F105 D0:F104 vdd vdd PSVTGP L=0.06u W=0.82u ad=0.0861p as=0.0898116p lpe=3 ngcon=1 nrd=0.292683 nrs=0.292683 pd=0.21u po2act=0.464914 ps=0.365404u sca=2.07813 scb=0.000807962 scc=4.50361e-06
MMMP15 net5:F141 D1:F140 vdd vdd PSVTGP L=0.06u W=0.82u ad=0.082p as=0.082p lpe=3 ngcon=1 nrd=0.268293 nrs=0.268293 pd=0.2u po2act=1.86096 ps=0.2u sca=2.07299 scb=0.000807962 scc=4.50361e-06
MMMP15@2 net5:F143 D1:F144 vdd vdd PSVTGP AD=0.082p AS=0.082p L=0.06u NRD=0.268293 NRS=0.268293 PD=0.2u PS=0.2u W=0.82u lpe=3 ngcon=1 po2act=1.86096 sca=2.07344 scb=0.000807962 scc=4.50361e-06
MMMP15@3 net5:F149 D1:F148 vdd vdd PSVTGP L=0.06u W=0.82u ad=0.082p as=0.0855875p lpe=3 ngcon=1 nrd=0.268293 nrs=0.268293 pd=0.2u po2act=1.78866 ps=0.290417u sca=2.07404 scb=0.000807962 scc=4.50361e-06
MMMP16 net8:F117 S0:F116 net16:F115 vdd PSVTGP L=0.06u W=0.82u ad=0.1476p as=0.082p lpe=3 ngcon=1 nrd=0.292683 nrs=0.268293 pd=1.18u po2act=0.342674 ps=0.2u sca=2.07323 scb=0.000807962 scc=4.50361e-06
MMMP16@2 net8:F119 S0:F120 net16:F121 vdd PSVTGP AD=0.082p AS=0.082p L=0.06u NRD=0.268293 NRS=0.268293 PD=0.2u PS=0.2u W=0.82u lpe=3 ngcon=1 po2act=0.776471 sca=2.07284 scb=0.000807962 scc=4.50361e-06
MMMP16@3 net8:F125 S0:F124 net16:F123 vdd PSVTGP L=0.06u W=0.82u ad=0.082p as=0.082p lpe=3 ngcon=1 nrd=0.268293 nrs=0.268293 pd=0.2u po2act=1.13797 ps=0.2u sca=2.0726 scb=0.000807962 scc=4.50361e-06
MMMP17 net5:F127 net20:F128 net16:F129 vdd PSVTGP AD=0.082p AS=0.082p L=0.06u NRD=0.268293 NRS=0.268293 PD=0.2u PS=0.2u W=0.82u lpe=3 ngcon=1 po2act=1.42717 sca=2.07249 scb=0.000807962 scc=4.50361e-06
MMMP17@2 net5:F133 net20:F132 net16:F131 vdd PSVTGP L=0.06u W=0.82u ad=0.082p as=0.082p lpe=3 ngcon=1 nrd=0.268293 nrs=0.268293 pd=0.2u po2act=1.64406 ps=0.2u sca=2.07252 scb=0.000807962 scc=4.50361e-06
MMMP17@3 net5:F135 net20:F136 net16:F137 vdd PSVTGP AD=0.082p AS=0.082p L=0.06u NRD=0.268293 NRS=0.268293 PD=0.2u PS=0.2u W=0.82u lpe=3 ngcon=1 po2act=1.78866 sca=2.07268 scb=0.000807962 scc=4.50361e-06
MMMP18 net20:F107 S0:F108 vdd vdd PSVTGP AD=0.075625p AS=0.0662634p L=0.06u NRD=0.421488 NRS=0.297521 PD=0.25u PS=0.269596u W=0.605u lpe=3 ngcon=1 po2act=0.655541 sca=2.41977 scb=0.00109035 scc=6.10399e-06
MMMP18@2 net20:F113 S0:F112 vdd vdd PSVTGP L=0.06u W=0.605u ad=0.075625p as=0.1089p lpe=3 ngcon=1 nrd=0.371901 nrs=0.297521 pd=0.25u po2act=0.316216 ps=0.965u sca=2.41814 scb=0.00109035 scc=6.10399e-06
R1 net8:F97 net8:F125 361.767
R10 net8:F105 net8:F99 0.001
R100 net20:F48 net20:F40 273.798
R101 net20:F48 net20:F31 350.683
R102 net20:F44 net20:F40 123.499
R103 net20:F44 net20:F31 400.405
R104 net20:F40 net20:F31 780.791
R105 net20:F31 net20:F37 0.001
R106 Z Z:F6 0.001
R107 Z:F6 Z:F167 19.359
R108 Z:F6 Z:F165 19.2285
R109 Z:F6 Z:F157 19.4546
R11 net8:F105 net8:F49 336.989
R110 Z:F6 Z:F91 19.1679
R111 Z:F6 Z:F89 19.2418
R112 Z:F6 Z:F81 19.4424
R113 Z:F157 Z:F167 2288.46
R114 Z:F157 Z:F165 2273.03
R115 Z:F157 Z:F151 0.001
R116 Z:F165 Z:F167 2261.87
R117 Z:F165 Z:F159 0.001
R118 Z:F81 Z:F89 1108.89
R119 Z:F81 Z:F75 0.001
R12 net8:F105 net8:F41 335.794
R120 Z:F89 Z:F83 0.001
R121 vdd vdd 0.001
R122 vdd vdd 42.8685
R123 vdd vdd 42.7242
R124 vdd vdd 42.9648
R125 vdd vdd 42.96
R126 vdd vdd 39.6854
R127 vdd vdd 39.5528
R128 vdd vdd 37.548
R129 vdd vdd 1423.91
R13 net8:F105 net8:F29 288.802
R130 vdd vdd 1419.12
R131 vdd vdd 1427.11
R132 vdd vdd 0.001
R133 vdd vdd 4645.8
R134 vdd vdd 4563.69
R135 vdd vdd 1424.07
R136 vdd vdd 1419.28
R137 vdd vdd 0.001
R138 vdd vdd 3539.49
R139 vdd vdd 4564.2
R14 net8:F105 net8:F21 294.721
R140 vdd vdd 1416.1
R141 vdd vdd 0.001
R142 vdd vdd 4620.3
R143 vdd vdd 4538.64
R144 vdd vdd 0.001
R145 vdd vdd 4635.9
R146 vdd vdd 4553.97
R147 vdd vdd 0.001
R148 vdd vdd 0.001
R149 vdd vdd 0.001
R15 net8:F117 net8:F125 256.888
R150 vdd vdd 0.001
R151 vdd vdd 0.001
R152 vdd vdd 0.001
R153 vdd vdd 0.001
R154 vdd vdd 0.001
R155 vdd vdd 0.001
R156 vdd vdd 0.001
R157 vdd vdd 0.001
R158 vdd vdd 0.001
R159 vdd vdd 0.001
R16 net8:F117 net8:F49 283.492
R160 vdd vdd 0.001
R161 vdd vdd 0.001
R162 vdd vdd 0.001
R163 vdd vdd 0.001
R164 vdd vdd 0.001
R165 vdd vdd 0.001
R166 vdd vdd 0.001
R167 vdd vdd 0.001
R168 vdd vdd 0.001
R169 vdd vdd 37.6272
R17 net8:F117 net8:F41 281.323
R170 D1 D1:F4 0.001
R171 D1:F68 D1:F148 634.612
R172 D1:F68 D1:F144 359.756
R173 D1:F68 D1:F140 680.421
R174 D1:F68 D1:F72 1035.42
R175 D1:F68 D1:F64 1110.16
R176 D1:F68 D1:F4 285.071
R177 D1:F148 D1:F144 388.956
R178 D1:F148 D1:F140 735.648
R179 D1:F148 D1:F72 229.455
R18 net8:F117 net8:F29 326.673
R180 D1:F148 D1:F64 1200.27
R181 D1:F148 D1:F4 308.209
R182 D1:F140 D1:F144 417.032
R183 D1:F140 D1:F72 1200.27
R184 D1:F140 D1:F64 219.913
R185 D1:F140 D1:F4 330.457
R186 D1:F144 D1:F72 634.612
R187 D1:F144 D1:F64 680.421
R188 D1:F144 D1:F4 174.721
R189 D1:F64 D1:F72 1958.33
R19 net8:F117 net8:F21 333.368
R190 D1:F64 D1:F4 539.167
R191 D1:F4 D1:F72 502.868
R192 gnd gnd 0.001
R193 gnd gnd 0.0256454
R194 gnd gnd 37.6237
R195 gnd gnd 0.001
R196 gnd gnd 0.001
R197 gnd gnd 0.001
R198 gnd gnd 0.001
R199 gnd gnd 0.001
R2 net8:F97 net8:F117 355.432
R20 net8:F125 net8:F119 0.001
R200 gnd gnd 0.001
R201 gnd gnd 0.001
R202 gnd gnd 0.001
R203 gnd gnd 0.001
R204 gnd gnd 0.001
R205 gnd gnd 0.001
R206 gnd gnd 0.001
R207 gnd gnd 0.001
R208 gnd gnd 0.001
R209 gnd gnd 0.001
R21 net8:F125 net8:F49 288.544
R210 gnd gnd 0.001
R211 gnd gnd 0.001
R212 gnd gnd 0.001
R213 S0 S0:F5 0.001
R214 S0:F5 S0:F124 1793.61
R215 S0:F5 S0:F120 876.875
R216 S0:F5 S0:F116 342.99
R217 S0:F5 S0:F112 78.731
R218 S0:F5 S0:F108 96.5919
R219 S0:F5 S0:F36 437.315
R22 net8:F125 net8:F41 286.337
R220 S0:F5 S0:F32 298.557
R221 S0:F124 S0:F120 115.74
R222 S0:F124 S0:F116 285.477
R223 S0:F124 S0:F112 1959.68
R224 S0:F124 S0:F108 5269.77
R225 S0:F124 S0:F36 10885.1
R226 S0:F124 S0:F32 16288.4
R227 S0:F56 S0:F60 207.605
R228 S0:F56 S0:F52 222.411
R229 S0:F56 S0:F36 1542.68
R23 net8:F125 net8:F29 332.494
R230 S0:F60 S0:F52 325.989
R231 S0:F60 S0:F36 2261.11
R232 S0:F52 S0:F36 839.138
R233 S0:F36 S0:F120 5321.63
R234 S0:F36 S0:F116 2081.55
R235 S0:F36 S0:F112 477.807
R236 S0:F36 S0:F108 1284.87
R237 S0:F36 S0:F32 3971.41
R238 S0:F116 S0:F120 139.566
R239 S0:F116 S0:F112 374.748
R24 net8:F125 net8:F21 339.309
R240 S0:F116 S0:F108 1007.73
R241 S0:F116 S0:F32 3114.81
R242 S0:F120 S0:F112 958.067
R243 S0:F120 S0:F108 2576.33
R244 S0:F120 S0:F32 7963.2
R245 S0:F108 S0:F112 231.318
R246 S0:F108 S0:F32 211.534
R247 S0:F112 S0:F32 714.983
R248 gnd gnd 0.001
R249 gnd gnd 4845.63
R25 net8:F21 net8:F49 320.778
R250 gnd gnd 4821.87
R251 gnd gnd 4579.56
R252 gnd gnd 5.68181
R253 gnd gnd 10.8616
R254 gnd gnd 10.2111
R255 gnd gnd 1832.12
R256 gnd gnd 1836.03
R257 gnd gnd 1837.29
R258 gnd gnd 0.001
R259 gnd gnd 4472.12
R26 net8:F21 net8:F41 319.641
R260 gnd gnd 4489.55
R261 gnd gnd 41.9708
R262 gnd gnd 1846.27
R263 gnd gnd 1850.21
R264 gnd gnd 0.001
R265 gnd gnd 4506.67
R266 gnd gnd 4524.24
R267 gnd gnd 42.2951
R268 gnd gnd 1845
R269 gnd gnd 0.001
R27 net8:F21 net8:F29 274.91
R270 gnd gnd 4503.58
R271 gnd gnd 4521.13
R272 gnd gnd 42.266
R273 gnd gnd 0.001
R274 gnd gnd 4493.99
R275 gnd gnd 4511.5
R276 gnd gnd 42.176
R277 gnd gnd 39.8814
R278 gnd gnd 40.0368
R279 gnd gnd 37.7185
R28 net8:F29 net8:F49 314.336
R280 gnd gnd 0.001
R281 gnd gnd 4266.04
R282 gnd gnd 0.001
R283 net16:375 net16:F168 5289.12
R284 net16:375 net16:F164 1880.83
R285 net16:375 net16:F160 544.14
R286 net16:375 net16:F156 174.94
R287 net16:375 net16:F152 147.701
R288 net16:375 net16:F137 37.5
R289 net16:375 net16:F129 38.9262
R29 net8:F29 net8:F41 313.222
R290 net16:375 net16:F121 39.6735
R291 net16:375 net16:F92 4848.36
R292 net16:375 net16:F88 1724.09
R293 net16:375 net16:F84 498.795
R294 net16:375 net16:F80 160.362
R295 net16:375 net16:F76 135.393
R296 net16:375 net16:F61 54.911
R297 net16:375 net16:F53 56.8746
R298 net16:375 net16:F45 57.9005
R299 net16:F160 net16:F168 1128.52
R3 net8:F97 net8:F105 245.576
R30 net8:F29 net8:F23 0.001
R300 net16:F160 net16:F164 401.307
R301 net16:F160 net16:F156 426.444
R302 net16:F160 net16:F152 1422.52
R303 net16:F160 net16:F92 1034.48
R304 net16:F160 net16:F88 371.735
R305 net16:F160 net16:F84 107.546
R306 net16:F160 net16:F80 390.907
R307 net16:F160 net16:F76 1303.97
R308 net16:F160 net16:F61 9359.96
R309 net16:F160 net16:F53 9694.66
R31 net8:F41 net8:F49 301.593
R310 net16:F160 net16:F45 9869.54
R311 net16:F164 net16:F168 310.005
R312 net16:F164 net16:F156 1474.01
R313 net16:F164 net16:F152 4916.96
R314 net16:F164 net16:F92 284.171
R315 net16:F164 net16:F88 101.052
R316 net16:F164 net16:F84 371.735
R317 net16:F164 net16:F80 1351.18
R318 net16:F164 net16:F76 4507.21
R319 net16:F168 net16:F156 4145.1
R32 net8:F49 net8:F43 0.001
R320 net16:F168 net16:F152 13827.1
R321 net16:F168 net16:F92 80.268
R322 net16:F168 net16:F88 284.171
R323 net16:F168 net16:F84 1045.36
R324 net16:F168 net16:F80 3799.67
R325 net16:F168 net16:F76 12674.8
R326 net16:F137 net16:F131 0.001
R327 net16:F152 net16:F156 457.338
R328 net16:F152 net16:F92 12674.8
R329 net16:F152 net16:F88 4507.21
R33 D0 D0:F3 0.001
R330 net16:F152 net16:F84 1303.97
R331 net16:F152 net16:F80 419.227
R332 net16:F152 net16:F76 101.962
R333 net16:F152 net16:F61 2540.67
R334 net16:F152 net16:F53 2631.52
R335 net16:F152 net16:F45 2678.99
R336 net16:F156 net16:F92 3799.67
R337 net16:F156 net16:F88 1351.18
R338 net16:F156 net16:F84 390.907
R339 net16:F156 net16:F80 125.676
R34 D0:F100 D0:F104 2073.02
R340 net16:F156 net16:F76 419.227
R341 net16:F156 net16:F61 3009.22
R342 net16:F156 net16:F53 3116.82
R343 net16:F156 net16:F45 3173.05
R344 net16:F84 net16:F92 958.251
R345 net16:F84 net16:F88 340.757
R346 net16:F84 net16:F80 358.332
R347 net16:F84 net16:F76 1195.31
R348 net16:F84 net16:F61 8579.96
R349 net16:F84 net16:F53 8886.77
R35 D0:F100 D0:F96 2603.96
R350 net16:F84 net16:F45 9047.08
R351 net16:F88 net16:F92 260.49
R352 net16:F88 net16:F80 1238.58
R353 net16:F88 net16:F76 4131.61
R354 net16:F88 net16:F61 13872.3
R355 net16:F88 net16:F53 14368.4
R356 net16:F88 net16:F45 14627.6
R357 net16:F92 net16:F80 3483.04
R358 net16:F92 net16:F76 11618.6
R359 net16:F76 net16:F80 384.291
R36 D0:F100 D0:F28 584.698
R360 net16:F76 net16:F61 2328.95
R361 net16:F76 net16:F53 2412.22
R362 net16:F76 net16:F45 2455.74
R363 net16:F80 net16:F61 2758.45
R364 net16:F80 net16:F53 2857.09
R365 net16:F80 net16:F45 2908.63
R366 net16:F61 net16:F55 0.001
R367 net16:F61 net16:F53 455.445
R368 net16:F61 net16:F45 463.661
R369 net16:F121 net16:F129 2066.67
R37 D0:F100 D0:F24 268.201
R370 net16:F121 net16:F115 0.001
R371 net16:F129 net16:F123 0.001
R372 net16:F45 net16:F53 393.935
R373 net16:F45 net16:F39 0.001
R374 net16:F53 net16:F47 0.001
R38 D0:F100 D0:F20 734.451
R39 D0:F100 D0:F3 650.209
R4 net8:F97 net8:F49 342.009
R40 D0:F104 D0:F96 5676.82
R41 D0:F104 D0:F28 195.507
R42 D0:F104 D0:F24 584.698
R43 D0:F104 D0:F20 1601.16
R44 D0:F104 D0:F3 1417.5
R45 D0:F96 D0:F28 1601.16
R46 D0:F96 D0:F24 734.451
R47 D0:F96 D0:F20 221.193
R48 D0:F96 D0:F3 522.457
R49 D0:F3 D0:F28 399.808
R5 net8:F97 net8:F41 340.797
R50 D0:F3 D0:F24 183.392
R51 D0:F3 D0:F20 147.36
R52 D0:F20 D0:F28 451.608
R53 D0:F20 D0:F24 207.153
R54 D0:F24 D0:F28 164.915
R55 net5:F133 net5:F149 221.573
R56 net5:F133 net5:F141 218.163
R57 net5:F133 net5:F127 0.001
R58 net5:F133 net5:F73 239.115
R59 net5:F133 net5:F65 235.112
R6 net8:F97 net8:F29 293.105
R60 net5:F133 net5:F57 239.484
R61 net5:F141 net5:F149 217.81
R62 net5:F141 net5:F135 0.001
R63 net5:F141 net5:F73 235.054
R64 net5:F141 net5:F65 231.119
R65 net5:F141 net5:F57 235.418
R66 net5:F149 net5:F143 0.001
R67 net5:F149 net5:F73 238.728
R68 net5:F149 net5:F65 234.732
R69 net5:F149 net5:F57 239.097
R7 net8:F97 net8:F21 299.112
R70 net5:F57 net5:F73 222.152
R71 net5:F57 net5:F65 218.433
R72 net5:F57 net5:F51 0.001
R73 net5:F65 net5:F73 218.096
R74 net5:F65 net5:F59 0.001
R75 net5:F73 net5:F67 0.001
R76 net20:F107 net20:F136 685.798
R77 net20:F107 net20:F132 380.999
R78 net20:F107 net20:F128 331.324
R79 net20:F107 net20:F113 0.001
R8 net8:F105 net8:F125 356.456
R80 net20:F107 net20:F48 332.912
R81 net20:F107 net20:F44 380.115
R82 net20:F107 net20:F40 741.224
R83 net20:F107 net20:F31 163.201
R84 net20:F132 net20:F136 116.612
R85 net20:F132 net20:F128 141.2
R86 net20:F132 net20:F48 613.408
R87 net20:F132 net20:F44 700.382
R88 net20:F132 net20:F40 1365.74
R89 net20:F132 net20:F31 401.337
R9 net8:F105 net8:F117 350.215
R90 net20:F136 net20:F128 254.16
R91 net20:F136 net20:F48 1104.13
R92 net20:F136 net20:F44 1260.69
R93 net20:F136 net20:F40 2458.34
R94 net20:F136 net20:F31 722.406
R95 net20:F128 net20:F48 533.431
R96 net20:F128 net20:F44 609.066
R97 net20:F128 net20:F40 1187.68
R98 net20:F128 net20:F31 349.01
R99 net20:F48 net20:F44 140.409
.ENDS HS65_GS_MUX21X44


.SUBCKT HS65_GS_NAND2X7 Z B A gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:19 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=2.044 PJ=5.72
MMM64 net247:F15 A:F16 gnd gnd NSVTGP AD=0.0624p AS=0.1521p L=0.06u NRD=0.102564 NRS=0.307692 PD=0.16u PS=1.17u W=0.78u lpe=3 ngcon=1 po2act=0.265328 sca=6.99475 scb=0.00671895 scc=0.000548722
MMM65 Z:F23 A:F24 vdd vdd PSVTGP AD=0.11p AS=0.1925p L=0.06u NRD=0.125 NRS=0.25 PD=0.2u PS=1.45u W=1.1u lpe=3 ngcon=1 po2act=0.24959 sca=5.22747 scb=0.00477169 scc=0.000389094
MMM66 Z:F29 B:F28 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.1925p lpe=3 ngcon=1 nrd=0.125 nrs=0.25 pd=0.2u po2act=0.24959 ps=1.45u sca=5.22747 scb=0.00477169 scc=0.000389094
MMM67 Z:F19 B:F20 net247:F21 gnd NSVTGP AD=0.1521p AS=0.0624p L=0.06u NRD=0.307692 NRS=0.102564 PD=1.17u PS=0.16u W=0.78u lpe=3 ngcon=1 po2act=0.265328 sca=6.99475 scb=0.00671895 scc=0.000548722
R1 net247:F15 net247:F21 0.001
R10 B:F28 B:F4 105.86
R11 B:F4 B:F20 92.5077
R12 A A:F3 0.001
R13 A:F24 A:F3 106.071
R14 A:F24 A:F16 62.2215
R15 A:F3 A:F16 92.6927
R16 vdd vdd 0.001
R17 vdd vdd 0.001
R18 vdd vdd 0.001
R19 vdd vdd 37.6252
R2 gnd gnd 0.001
R20 vdd vdd 0.001
R21 vdd vdd 37.6266
R22 vdd vdd 37.5
R23 gnd gnd 0.001
R24 gnd gnd 0.0256454
R25 gnd gnd 37.6237
R26 gnd gnd 0.001
R3 gnd gnd 37.5194
R4 Z Z:F5 0.001
R5 Z:F23 Z:F29 0.001
R6 Z:F23 Z:F5 20.2347
R7 Z:F5 Z:F19 37.5
R8 B B:F4 0.001
R9 B:F28 B:F20 62.2604
.ENDS HS65_GS_NAND2X7


.SUBCKT HS65_GS_NOR2AX3 Z B A gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:21 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=2.336 PJ=6.12
MMM29 net091:F18 A:F17 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.07515p as=0.0213846p lpe=3 ngcon=1 nrd=3.08333 nrs=0.275 pd=1.39u po2act=0.244444 ps=0.2u sca=17.6177 scb=0.0199621 scc=0.00206349
MMM31 net091:F30 A:F29 vdd vdd PSVTGP L=0.06u W=0.29u ad=0.04785p as=0.0675976p lpe=3 ngcon=1 nrd=0.189655 nrs=2.15712 pd=0.62u po2act=0.157333 ps=0.776786u sca=9.72382 scb=0.0116961 scc=0.00066791
MMM64 Z:F26 B:F25 gnd gnd NSVTGP L=0.06u W=0.32u ad=0.032p as=0.10915p lpe=3 ngcon=1 nrd=0.34375 nrs=2.27083 pd=0.2u po2act=0.221307 ps=1.81u sca=13.2913 scb=0.0149125 scc=0.0013319
MMM65 net0156:F32 net091:F33 vdd vdd PSVTGP AD=0.0385p AS=0.128202p L=0.06u NRD=0.127273 NRS=0.105195 PD=0.14u PS=1.47321u W=0.55u lpe=3 ngcon=1 po2act=0.224015 sca=1.86996 scb=0.000422129 scc=6.91737e-07
MMM66 Z:F36 B:F37 net0156:F38 vdd PSVTGP AD=0.09075p AS=0.0385p L=0.06u NRD=0.3 NRS=0.127273 PD=0.88u PS=0.14u W=0.55u lpe=3 ngcon=1 po2act=0.227882 sca=1.87015 scb=0.000422129 scc=6.91737e-07
MMM67 Z:F20 net091:F21 gnd gnd NSVTGP AD=0.032p AS=0.0342154p L=0.06u NRD=0.34375 NRS=0.34375 PD=0.2u PS=0.32u W=0.32u lpe=3 ngcon=1 po2act=0.289477 sca=13.2912 scb=0.0149125 scc=0.0013319
R1 gnd gnd 0.001
R10 Z:F5 Z:F20 37.9229
R11 Z:F20 Z:F26 0.001
R12 B B:F4 0.001
R13 B:F37 B:F4 65.6278
R14 B:F37 B:F25 199.893
R15 B:F4 B:F25 358.112
R16 net091:F33 net091:F30 972.002
R17 net091:F33 net091:F21 210.581
R18 net091:F33 net091:F18 982.665
R19 net091:F30 net091:F21 183.625
R2 gnd gnd 37.7139
R20 net091:F30 net091:F18 100.752
R21 net091:F21 net091:F18 185.639
R22 net0156:F32 net0156:F38 0.001
R23 vdd vdd 0.001
R24 vdd vdd 0.001
R25 vdd vdd 0.001
R26 vdd vdd 0.001
R27 vdd vdd 37.6252
R28 vdd vdd 0.001
R29 vdd vdd 18.7759
R3 gnd gnd 38.2936
R30 vdd vdd 0.001
R31 gnd gnd 0.001
R32 gnd gnd 0.001
R33 gnd gnd 0.001
R34 gnd gnd 0.0256454
R35 gnd gnd 37.6237
R4 gnd gnd 0.001
R5 A A:F3 0.001
R6 A:F3 A:F29 48.6273
R7 A:F29 A:F17 78.1521
R8 Z Z:F5 0.001
R9 Z:F36 Z:F5 39.5899
.ENDS HS65_GS_NOR2AX3


.SUBCKT HS65_GS_NOR2X6 Z B A gnd gnd vdd vdd
*modified
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:22 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=2.044 PJ=5.72
MMM64 Z:F21 B:F20 gnd gnd NSVTGP L=0.06u W=0.63u ad=0.063p as=0.11025p lpe=3 ngcon=1 nrd=0.130952 nrs=0.261905 pd=0.2u po2act=0.24959 ps=0.98u sca=4.02706 scb=0.00326609 scc=7.50079e-05
MMM65 net0156:F23 A:F24 vdd vdd PSVTGP AD=0.0935p AS=0.209p L=0.06u NRD=0.0772727 NRS=0.295455 PD=0.17u PS=1.48u W=1.1u lpe=3 ngcon=1 po2act=0.261639 sca=5.22746 scb=0.00477169 scc=0.000389094
MMM66 Z:F27 B:F28 net0156:F29 vdd PSVTGP AD=0.209p AS=0.0935p L=0.06u NRD=0.272727 NRS=0.0772727 PD=1.48u PS=0.17u W=1.1u lpe=3 ngcon=1 po2act=0.261639 sca=5.22746 scb=0.00477169 scc=0.000389094
MMM67 Z:F15 A:F16 gnd gnd NSVTGP AD=0.063p AS=0.11025p L=0.06u NRD=0.130952 NRS=0.261905 PD=0.2u PS=0.98u W=0.63u lpe=3 ngcon=1 po2act=0.24959 sca=4.02706 scb=0.00326609 scc=7.50079e-05
R1 gnd gnd 0.001
R10 B:F28 B:F4 83.3323
R11 B:F4 B:F20 171.022
R12 A A:F3 0.001
R13 A:F24 A:F16 124.069
R14 A:F24 A:F3 83.3341
R15 A:F3 A:F16 171.026
R16 net0156:F23 net0156:F29 0.001
R17 vdd vdd 0.001
R18 vdd vdd 0.001
R19 vdd vdd 0.001
R2 gnd gnd 37.5
R20 vdd vdd 37.6252
R21 vdd vdd 0.001
R22 vdd vdd 37.5
R23 gnd gnd 0.001
R24 gnd gnd 0.0256454
R25 gnd gnd 37.6237
R26 gnd gnd 0.001
R3 gnd gnd 37.6187
R4 Z Z:F5 0.001
R5 Z:F27 Z:F5 39.0608
R6 Z:F5 Z:F15 18.8987
R7 Z:F15 Z:F21 0.001
R8 B B:F4 0.001
R9 B:F28 B:F20 124.071
.ENDS HS65_GS_NOR2X6


.SUBCKT HS65_GS_NOR4ABX2 Z D C B A gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:23 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=2.92 PJ=6.92
MMM0 net013:F48 net042:F49 vdd vdd PSVTGP AD=0.028275p AS=0.0922626p L=0.06u NRD=0.149425 NRS=0.321839 PD=0.13u PS=1.1529u W=0.435u lpe=3 ngcon=1 po2act=0.264026 sca=1.3278 scb=6.51395e-05 scc=1.00045e-08
MMM1 Z:F32 net042:F33 gnd gnd NSVTGP AD=0.0509833p AS=0.0255p L=0.06u NRD=0.275 NRS=0.325 PD=0.62u PS=0.255u W=0.2u lpe=3 ngcon=1 po2act=0.275305 sca=17.6157 scb=0.0199621 scc=0.00206349
MMM2 Z:F38 C:F37 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0509833p as=0.035p lpe=3 ngcon=1 nrd=1.99753 nrs=0.275 pd=0.62u po2act=0.169853 ps=0.55u sca=3.30122 scb=0.0017987 scc=7.29807e-06
MMM24 net042:F40 B:F41 vdd vdd PSVTGP AD=0.028p AS=0.138125p L=0.06u NRD=0.196429 NRS=3.71296 PD=0.2u PS=2.34u W=0.28u lpe=3 ngcon=1 po2act=0.208534 sca=9.91523 scb=0.0119886 scc=0.000690876
MMM25 net042:F46 A:F45 vdd vdd PSVTGP L=0.06u W=0.28u ad=0.028p as=0.0593874p lpe=3 ngcon=1 nrd=0.196429 nrs=3.05061 pd=0.2u po2act=0.216505 ps=0.742098u sca=9.91471 scb=0.0119886 scc=0.000690876
MMM26 net042:F22 B:F21 net45:F20 gnd NSVTGP L=0.06u W=0.2u ad=0.0733p as=0.013p lpe=3 ngcon=1 nrd=2.68148 nrs=0.325 pd=1.37u po2act=0.232195 ps=0.13u sca=17.6161 scb=0.0199621 scc=0.00206349
MMM27 net45:F26 A:F25 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.013p as=0.0255p lpe=3 ngcon=1 nrd=0.325 nrs=0.5 pd=0.13u po2act=0.39439 ps=0.255u sca=17.6159 scb=0.0199621 scc=0.00206349
MMM3 Z:F28 D:F29 gnd gnd NSVTGP AD=0.0509833p AS=0.038p L=0.06u NRD=7.045 NRS=0.325 PD=0.62u PS=0.58u W=0.2u lpe=3 ngcon=1 po2act=0.239806 sca=1.88934 scb=0.000214041 scc=7.20983e-08
MMM4 net041:F52 C:F53 net013:F54 vdd PSVTGP AD=0.028275p AS=0.028275p L=0.06u NRD=0.149425 NRS=0.149425 PD=0.13u PS=0.13u W=0.435u lpe=3 ngcon=1 po2act=0.361092 sca=1.32798 scb=6.51395e-05 scc=1.00045e-08
MMM5 Z:F56 D:F57 net041:F58 vdd PSVTGP AD=0.071775p AS=0.028275p L=0.06u NRD=0.252874 NRS=0.149425 PD=0.765u PS=0.13u W=0.435u lpe=3 ngcon=1 po2act=0.254736 sca=1.32837 scb=6.51395e-05 scc=1.00045e-08
R1 net45:F20 net45:F26 0.001
R10 B B:F4 0.001
R11 B:F4 B:F41 137.723
R12 B:F4 B:F21 86.6752
R13 B:F41 B:F21 93.3748
R14 A A:F3 0.001
R15 A:F3 A:F45 116.089
R16 A:F45 A:F25 110
R17 Z Z:F7 0.001
R18 Z:F56 Z:F7 37.8073
R19 Z:F7 Z:F32 39.1472
R2 gnd gnd 0.001
R20 Z:F32 Z:F38 0.001
R21 Z:F32 Z:F28 0.001
R22 net041:F52 net041:F58 0.001
R23 D D:F6 0.001
R24 D:F57 D:F29 3438.44
R25 D:F57 D:F6 322.81
R26 D:F6 D:F29 495.694
R27 C C:F5 0.001
R28 C:F53 C:F37 715.752
R29 C:F53 C:F5 132.908
R3 gnd gnd 38.1438
R30 C:F5 C:F37 337.091
R31 net013:F48 net013:F54 0.001
R32 net042:F49 net042:F46 920.659
R33 net042:F49 net042:F33 341.331
R34 net042:F49 net042:F22 944.39
R35 net042:F46 net042:F40 0.001
R36 net042:F46 net042:F33 222.056
R37 net042:F46 net042:F22 96.9979
R38 net042:F33 net042:F22 227.78
R39 vdd vdd 0.001
R4 gnd gnd 37.8537
R40 vdd vdd 0.001
R41 vdd vdd 0.001
R42 vdd vdd 0.001
R43 vdd vdd 0.001
R44 vdd vdd 0.001
R45 vdd vdd 37.6252
R46 vdd vdd 0.001
R47 vdd vdd 37.6254
R48 vdd vdd 37.534
R49 vdd vdd 0.001
R5 gnd gnd 38.5745
R50 gnd gnd 0.001
R51 gnd gnd 0.001
R52 gnd gnd 0.001
R53 gnd gnd 0.001
R54 gnd gnd 0.001
R55 gnd gnd 0.0256454
R56 gnd gnd 37.6237
R6 gnd gnd 13072.2
R7 gnd gnd 0.001
R8 gnd gnd 12972.7
R9 gnd gnd 12827.9
.ENDS HS65_GS_NOR4ABX2


.SUBCKT HS65_GS_OAI21X3 Z C B A gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:28 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=2.336 PJ=6.12
MMM43 Z:F33 B:F34 net0158:F35 vdd PSVTGP AD=0.056375p AS=0.039875p L=0.06u NRD=0.3 NRS=0.131818 PD=0.205u PS=0.145u W=0.55u lpe=3 ngcon=1 po2act=0.402778 sca=1.48303 scb=0.000143767 scc=6.83223e-08
MMM47 Z:F39 C:F38 vdd vdd PSVTGP L=0.06u W=0.55u ad=0.056375p as=0.0935p lpe=3 ngcon=1 nrd=0.327273 nrs=0.3 pd=0.205u po2act=0.268642 ps=0.89u sca=1.48322 scb=0.000143767 scc=6.83223e-08
MMM52 net0158:F29 A:F30 vdd vdd PSVTGP AD=0.039875p AS=0.0935p L=0.06u NRD=0.131818 NRS=0.3 PD=0.145u PS=0.89u W=0.55u lpe=3 ngcon=1 po2act=0.268642 sca=1.48322 scb=0.000143767 scc=6.83223e-08
MMM77 Z:F25 C:F26 net020:F27 gnd NSVTGP AD=0.0726p AS=0.0955016p L=0.06u NRD=0.25 NRS=0.493294 PD=0.77u PS=1.32u W=0.44u lpe=3 ngcon=1 po2act=0.173503 sca=3.04441 scb=0.00159776 scc=1.00392e-05
MMM78 net020:F21 B:F22 gnd gnd NSVTGP AD=0.0846492p AS=0.039p L=0.06u NRD=0.556536 NRS=0.282051 PD=1.17u PS=0.2u W=0.39u lpe=3 ngcon=1 po2act=0.233211 sca=11.6429 scb=0.0127786 scc=0.00109616
MMM79 net020:F19 A:F18 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0846492p as=0.039p lpe=3 ngcon=1 nrd=0.556536 nrs=0.282051 pd=1.17u po2act=0.213282 ps=0.2u sca=11.643 scb=0.0127786 scc=0.00109616
R1 gnd gnd 0.001
R10 C C:F5 0.001
R11 C:F38 C:F5 137.88
R12 C:F38 C:F26 875.29
R13 C:F5 C:F26 92.5803
R14 B B:F4 0.001
R15 B:F34 B:F22 298.821
R16 B:F34 B:F4 153.205
R17 B:F4 B:F22 146.977
R18 A A:F3 0.001
R19 A:F30 A:F18 351.148
R2 gnd gnd 38.0016
R20 A:F30 A:F3 431.941
R21 A:F3 A:F18 75.1171
R22 net0158:F29 net0158:F35 0.001
R23 vdd vdd 0.001
R24 vdd vdd 0.001
R25 vdd vdd 0.001
R26 vdd vdd 0.001
R27 vdd vdd 37.6252
R28 vdd vdd 0.001
R29 vdd vdd 37.6777
R3 gnd gnd 0.001
R30 vdd vdd 37.5
R31 gnd gnd 0.001
R32 gnd gnd 0.0256454
R33 gnd gnd 37.6237
R34 gnd gnd 0.001
R35 gnd gnd 0.001
R4 net020:F19 net020:F27 0.001
R5 net020:F19 net020:F21 0.001
R6 Z Z:F6 0.001
R7 Z:F33 Z:F39 0.001
R8 Z:F33 Z:F6 38.2069
R9 Z:F6 Z:F25 38.9009
.ENDS HS65_GS_OAI21X3


.SUBCKT HS65_GS_OAI21X37 Z C B A gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:28 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=8.176 PJ=14.12
MMM43 Z:F131 B:F130 net0158:F129 vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=2.33135 ps=0.2u sca=5.20642 scb=0.00477169 scc=0.000389094
MMM47 Z:F159 C:F158 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.209p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=0.364911 ps=1.48u sca=5.21364 scb=0.00477169 scc=0.000389094
MMM52 net0158:F89 A:F90 vdd vdd PSVTGP AD=0.11p AS=0.1925p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=1.45u W=1.1u lpe=3 ngcon=1 po2act=0.3372 sca=5.21396 scb=0.00477169 scc=0.000389094
MMM66 net0158:F95 A:F94 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=0.790909 ps=0.2u sca=5.21197 scb=0.00477169 scc=0.000389094
MMM67 Z:F109 B:F110 net0158:F111 vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=2.04065 sca=5.20728 scb=0.00477169 scc=0.000389094
MMM68 Z:F137 C:F138 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.125 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=2.05206 sca=5.20719 scb=0.00477169 scc=0.000389094
MMM69 net0158:F97 A:F98 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=1.18811 sca=5.21021 scb=0.00477169 scc=0.000389094
MMM70 Z:F115 B:F114 net0158:F113 vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=2.21181 ps=0.2u sca=5.20679 scb=0.00477169 scc=0.000389094
MMM71 Z:F143 C:F142 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.125 nrs=0.25 pd=0.2u po2act=1.82765 ps=0.2u sca=5.20783 scb=0.00477169 scc=0.000389094
MMM72 net0158:F103 A:F102 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=1.5288 ps=0.2u sca=5.2088 scb=0.00477169 scc=0.000389094
MMM73 Z:F117 B:F118 net0158:F119 vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=2.32646 sca=5.20646 scb=0.00477169 scc=0.000389094
MMM74 Z:F145 C:F146 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=1.54673 sca=5.20866 scb=0.00477169 scc=0.000389094
MMM75 net0158:F105 A:F106 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=1.81298 sca=5.20795 scb=0.00477169 scc=0.000389094
MMM76 Z:F123 B:F122 net0158:F121 vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=2.3846 ps=0.2u sca=5.20629 scb=0.00477169 scc=0.000389094
MMM77 Z:F87 C:F86 net020:F85 gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.1443p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=0.2u po2act=0.35568 ps=1.15u sca=6.98685 scb=0.00671895 scc=0.000548722
MMM78 net020:F59 B:F58 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=0.2u po2act=2.32798 ps=0.2u sca=6.98046 scb=0.00671895 scc=0.000548722
MMM79 net020:F19 A:F18 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.1365p as=0.078p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=1.13u po2act=0.337186 ps=0.2u sca=6.98706 scb=0.00671895 scc=0.000548722
MMM80 net020:F21 A:F22 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.282051 NRS=0.282051 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=0.790826 sca=6.98578 scb=0.00671895 scc=0.000548722
MMM81 net020:F37 B:F38 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.282051 NRS=0.282051 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=2.0397 sca=6.98175 scb=0.00671895 scc=0.000548722
MMM82 Z:F65 C:F66 net020:F67 gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.282051 NRS=0.282051 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=2.04731 sca=6.98163 scb=0.00671895 scc=0.000548722
MMM83 net020:F43 B:F42 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=0.2u po2act=2.21049 ps=0.2u sca=6.98096 scb=0.00671895 scc=0.000548722
MMM84 net020:F27 A:F26 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=0.2u po2act=1.1879 ps=0.2u sca=6.98462 scb=0.00671895 scc=0.000548722
MMM85 Z:F71 C:F70 net020:F69 gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=0.2u po2act=1.82212 ps=0.2u sca=6.98248 scb=0.00671895 scc=0.000548722
MMM86 Z:F73 C:F74 net020:F75 gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.282051 NRS=0.282051 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=1.54037 sca=6.98342 scb=0.00671895 scc=0.000548722
MMM87 net020:F29 A:F30 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.282051 NRS=0.282051 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=1.5284 sca=6.98357 scb=0.00671895 scc=0.000548722
MMM88 net020:F45 B:F46 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.282051 NRS=0.282051 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=2.32472 sca=6.98048 scb=0.00671895 scc=0.000548722
MMM89 net0158:F135 A:F134 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=2.21996 ps=0.2u sca=5.20672 scb=0.00477169 scc=0.000389094
MMM90 Z:F125 B:F126 net0158:F127 vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=2.38623 sca=5.20628 scb=0.00477169 scc=0.000389094
MMM91 Z:F151 C:F150 vdd vdd PSVTGP L=0.06u W=1.1u ad=0.11p as=0.11p lpe=3 ngcon=1 nrd=0.25 nrs=0.25 pd=0.2u po2act=1.2093 ps=0.2u sca=5.20996 scb=0.00477169 scc=0.000389094
MMM92 Z:F81 C:F82 net020:F83 gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.282051 NRS=0.282051 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=0.807144 sca=6.98559 scb=0.00671895 scc=0.000548722
MMM93 Z:F79 C:F78 net020:F77 gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=0.2u po2act=1.20204 ps=0.2u sca=6.98445 scb=0.00671895 scc=0.000548722
MMM94 net020:F35 A:F34 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=0.2u po2act=1.81233 ps=0.2u sca=6.98262 scb=0.00671895 scc=0.000548722
MMM95 net020:F61 A:F62 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.282051 NRS=0.282051 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=2.21593 sca=6.98085 scb=0.00671895 scc=0.000548722
MMM96 net020:F51 B:F50 gnd gnd NSVTGP L=0.06u W=0.78u ad=0.078p as=0.078p lpe=3 ngcon=1 nrd=0.282051 nrs=0.282051 pd=0.2u po2act=2.38237 ps=0.2u sca=6.98038 scb=0.00671895 scc=0.000548722
MMM97 net020:F53 B:F54 gnd gnd NSVTGP AD=0.078p AS=0.078p L=0.06u NRD=0.282051 NRS=0.282051 PD=0.2u PS=0.2u W=0.78u lpe=3 ngcon=1 po2act=2.38346 sca=6.98037 scb=0.00671895 scc=0.000548722
MMM98 Z:F153 C:F154 vdd vdd PSVTGP AD=0.11p AS=0.11p L=0.06u NRD=0.25 NRS=0.25 PD=0.2u PS=0.2u W=1.1u lpe=3 ngcon=1 po2act=0.815361 sca=5.21169 scb=0.00477169 scc=0.000389094
R1 net020:F53 net020:F85 387.399
R10 net020:F53 net020:F19 418.645
R100 Z:F65 Z:F71 0.001
R101 Z:F73 Z:F81 1538.22
R102 Z:F73 Z:F79 0.001
R103 Z:F81 Z:F87 0.001
R104 A A:F3 0.001
R105 A:F94 A:F106 4512.88
R106 A:F94 A:F102 1766.74
R107 A:F94 A:F98 392.617
R108 A:F94 A:F90 279.712
R109 A:F94 A:F34 4942.68
R11 net020:F61 net020:F85 354.811
R110 A:F94 A:F30 1935.01
R111 A:F94 A:F26 430.009
R112 A:F94 A:F22 116.809
R113 A:F94 A:F18 306.351
R114 A:F94 A:F3 144.106
R115 A:F134 A:F102 26315.2
R116 A:F134 A:F62 69.1296
R117 A:F134 A:F30 28821.4
R118 A:F134 A:F3 110.647
R119 A:F102 A:F106 271.927
R12 net020:F61 net020:F77 348.664
R120 A:F102 A:F98 404.212
R121 A:F102 A:F90 4633.59
R122 A:F102 A:F62 26315.2
R123 A:F102 A:F34 297.825
R124 A:F102 A:F30 116.595
R125 A:F102 A:F26 442.708
R126 A:F102 A:F22 1935.01
R127 A:F102 A:F18 5074.88
R128 A:F102 A:F3 147.373
R129 A:F62 A:F30 28821.4
R13 net020:F61 net020:F69 336.888
R130 A:F62 A:F3 110.647
R131 A:F106 A:F98 1032.5
R132 A:F106 A:F90 11835.8
R133 A:F106 A:F34 80.7863
R134 A:F106 A:F30 297.825
R135 A:F106 A:F26 1130.83
R136 A:F106 A:F22 4942.68
R137 A:F106 A:F18 12963
R138 A:F106 A:F3 372.271
R139 A:F3 A:F98 287.178
R14 net020:F61 net020:F67 0.001
R140 A:F3 A:F90 377.942
R141 A:F3 A:F34 407.726
R142 A:F3 A:F30 161.408
R143 A:F3 A:F26 314.528
R144 A:F3 A:F22 157.83
R145 A:F3 A:F18 413.936
R146 A:F22 A:F98 430.009
R147 A:F22 A:F90 306.351
R148 A:F22 A:F34 5413.41
R149 A:F22 A:F30 2119.29
R15 net020:F61 net020:F51 375.868
R150 A:F22 A:F26 470.963
R151 A:F22 A:F18 335.528
R152 A:F30 A:F98 442.708
R153 A:F30 A:F90 5074.88
R154 A:F30 A:F34 326.19
R155 A:F30 A:F26 484.871
R156 A:F30 A:F18 5558.2
R157 A:F90 A:F98 1029.71
R158 A:F90 A:F34 12963
R159 A:F90 A:F26 1127.77
R16 net020:F61 net020:F37 403.099
R160 A:F90 A:F18 80.0392
R161 A:F98 A:F34 1130.83
R162 A:F98 A:F26 98.3814
R163 A:F98 A:F18 1127.77
R164 A:F18 A:F34 14197.6
R165 A:F18 A:F26 1235.18
R166 A:F26 A:F34 1238.53
R167 vdd vdd 0.001
R168 vdd vdd 41.4731
R169 vdd vdd 41.6131
R17 net020:F61 net020:F29 423.858
R170 vdd vdd 41.1279
R171 vdd vdd 41.0586
R172 vdd vdd 38.9647
R173 vdd vdd 38.8657
R174 vdd vdd 37.5
R175 vdd vdd 2028.01
R176 vdd vdd 2034.86
R177 vdd vdd 2011.13
R178 vdd vdd 0.001
R179 vdd vdd 6070.64
R18 net020:F61 net020:F21 436.254
R180 vdd vdd 5999.87
R181 vdd vdd 2031.43
R182 vdd vdd 2038.29
R183 vdd vdd 0.001
R184 vdd vdd 6080.89
R185 vdd vdd 6010
R186 vdd vdd 2055.4
R187 vdd vdd 0.001
R188 vdd vdd 4594.42
R189 vdd vdd 6080.89
R19 net020:F61 net020:F19 446.495
R190 vdd vdd 6131.92
R191 vdd vdd 6060.43
R192 vdd vdd 0.001
R193 vdd vdd 0.001
R194 vdd vdd 0.001
R195 vdd vdd 0.001
R196 vdd vdd 0.001
R197 vdd vdd 0.001
R198 vdd vdd 0.001
R199 vdd vdd 0.001
R2 net020:F53 net020:F77 380.688
R20 net020:F69 net020:F85 322.043
R200 vdd vdd 0.001
R201 vdd vdd 0.001
R202 vdd vdd 0.001
R203 vdd vdd 0.001
R204 vdd vdd 0.001
R205 vdd vdd 0.001
R206 vdd vdd 0.001
R207 vdd vdd 0.001
R208 vdd vdd 0.001
R209 vdd vdd 0.001
R21 net020:F69 net020:F77 316.463
R210 vdd vdd 0.001
R211 vdd vdd 0.001
R212 vdd vdd 0.001
R213 vdd vdd 37.6252
R214 B B:F4 0.001
R215 B:F54 B:F130 291.751
R216 B:F54 B:F126 105.083
R217 B:F54 B:F122 443.087
R218 B:F54 B:F118 1743.01
R219 B:F54 B:F114 6561.45
R22 net020:F69 net020:F75 0.001
R220 B:F54 B:F58 319.537
R221 B:F54 B:F50 485.286
R222 B:F54 B:F46 1909.01
R223 B:F54 B:F42 7186.35
R224 B:F54 B:F4 236.536
R225 B:F38 B:F130 32270.9
R226 B:F38 B:F126 11623.3
R227 B:F38 B:F122 5431.37
R228 B:F38 B:F118 1529.33
R229 B:F38 B:F114 356.78
R23 net020:F69 net020:F51 395.19
R230 B:F38 B:F110 84.0092
R231 B:F38 B:F50 5948.64
R232 B:F38 B:F46 1674.98
R233 B:F38 B:F42 390.76
R234 B:F38 B:F4 202.894
R235 B:F42 B:F130 18217.2
R236 B:F42 B:F126 6561.45
R237 B:F42 B:F122 1602.71
R238 B:F42 B:F118 451.279
R239 B:F42 B:F114 105.28
R24 net020:F69 net020:F37 423.821
R240 B:F42 B:F110 356.78
R241 B:F42 B:F58 19952.2
R242 B:F42 B:F50 1755.35
R243 B:F42 B:F46 494.258
R244 B:F42 B:F4 184.491
R245 B:F46 B:F130 4839.29
R246 B:F46 B:F126 1743.01
R247 B:F46 B:F122 425.751
R248 B:F46 B:F118 119.88
R249 B:F46 B:F114 451.279
R25 net020:F69 net020:F29 445.647
R250 B:F46 B:F110 1529.33
R251 B:F46 B:F58 5300.18
R252 B:F46 B:F50 466.299
R253 B:F46 B:F4 136.085
R254 B:F50 B:F130 1230.19
R255 B:F50 B:F126 443.087
R256 B:F50 B:F122 106.671
R257 B:F50 B:F118 425.751
R258 B:F50 B:F114 1602.71
R259 B:F50 B:F110 5431.37
R26 net020:F69 net020:F21 458.68
R260 B:F50 B:F58 1347.35
R261 B:F50 B:F4 202.559
R262 B:F58 B:F130 77.7142
R263 B:F58 B:F126 291.751
R264 B:F58 B:F122 1230.19
R265 B:F58 B:F118 4839.29
R266 B:F58 B:F114 18217.2
R267 B:F58 B:F4 656.718
R268 B:F130 B:F126 266.381
R269 B:F130 B:F122 1123.21
R27 net020:F69 net020:F19 469.447
R270 B:F130 B:F118 4418.49
R271 B:F130 B:F114 16633.1
R272 B:F130 B:F110 29464.7
R273 B:F130 B:F4 599.612
R274 B:F122 B:F126 404.558
R275 B:F122 B:F118 388.729
R276 B:F122 B:F114 1463.34
R277 B:F122 B:F110 4959.08
R278 B:F122 B:F4 184.945
R279 B:F126 B:F118 1591.45
R28 net020:F77 net020:F85 290.133
R280 B:F126 B:F114 5990.89
R281 B:F126 B:F110 10612.6
R282 B:F126 B:F4 215.968
R283 B:F118 B:F114 412.038
R284 B:F118 B:F110 1396.34
R285 B:F118 B:F4 124.251
R286 B:F114 B:F110 325.756
R287 B:F114 B:F4 168.448
R288 B:F110 B:F4 185.251
R289 gnd gnd 0.001
R29 net020:F77 net020:F83 0.001
R290 gnd gnd 0.0256454
R291 gnd gnd 37.6237
R292 gnd gnd 0.001
R293 gnd gnd 0.001
R294 gnd gnd 0.001
R295 gnd gnd 0.001
R296 gnd gnd 0.001
R297 gnd gnd 0.001
R298 gnd gnd 0.001
R299 gnd gnd 0.001
R3 net020:F53 net020:F69 367.83
R30 net020:F77 net020:F51 409.004
R300 gnd gnd 0.001
R301 gnd gnd 0.001
R302 gnd gnd 0.001
R303 gnd gnd 0.001
R304 gnd gnd 0.001
R305 gnd gnd 0.001
R306 gnd gnd 0.001
R307 gnd gnd 0.001
R308 gnd gnd 0.001
R309 C C:F5 0.001
R31 net020:F77 net020:F37 438.636
R310 C:F5 C:F158 321.164
R311 C:F5 C:F154 129.188
R312 C:F5 C:F150 132.941
R313 C:F5 C:F146 428.382
R314 C:F5 C:F142 1470.8
R315 C:F5 C:F138 4105.88
R316 C:F5 C:F86 351.751
R317 C:F5 C:F82 141.491
R318 C:F5 C:F78 145.602
R319 C:F5 C:F74 407.983
R32 net020:F77 net020:F29 461.224
R320 C:F5 C:F70 1400.76
R321 C:F5 C:F66 3910.36
R322 C:F78 C:F158 1518.54
R323 C:F78 C:F154 610.831
R324 C:F78 C:F150 119.071
R325 C:F78 C:F146 383.688
R326 C:F78 C:F142 1317.35
R327 C:F78 C:F138 3677.5
R328 C:F78 C:F86 1663.17
R329 C:F78 C:F82 669.006
R33 net020:F77 net020:F21 474.714
R330 C:F78 C:F74 365.418
R331 C:F78 C:F70 1254.62
R332 C:F78 C:F66 3502.38
R333 C:F82 C:F158 288.327
R334 C:F82 C:F154 115.979
R335 C:F82 C:F150 610.832
R336 C:F82 C:F146 1968.32
R337 C:F82 C:F142 6757.98
R338 C:F82 C:F138 18865.5
R339 C:F82 C:F86 315.787
R34 net020:F77 net020:F19 485.857
R340 C:F82 C:F74 1874.59
R341 C:F82 C:F70 6436.17
R342 C:F82 C:F66 17967.2
R343 C:F146 C:F158 4467.78
R344 C:F146 C:F154 1797.16
R345 C:F146 C:F150 350.324
R346 C:F146 C:F142 340.98
R347 C:F146 C:F138 951.88
R348 C:F146 C:F86 4893.28
R349 C:F146 C:F74 94.5841
R35 net020:F85 net020:F51 416.215
R350 C:F146 C:F70 324.743
R351 C:F146 C:F66 906.552
R352 C:F150 C:F158 1386.5
R353 C:F150 C:F154 557.716
R354 C:F150 C:F142 1202.8
R355 C:F150 C:F138 3357.72
R356 C:F150 C:F86 1518.54
R357 C:F150 C:F74 333.642
R358 C:F150 C:F70 1145.52
R359 C:F150 C:F66 3197.83
R36 net020:F85 net020:F37 446.369
R360 C:F154 C:F158 263.255
R361 C:F154 C:F142 6170.33
R362 C:F154 C:F138 17225.1
R363 C:F154 C:F86 288.327
R364 C:F154 C:F74 1711.58
R365 C:F154 C:F70 5876.5
R366 C:F154 C:F66 16404.8
R367 C:F138 C:F142 264.578
R368 C:F138 C:F74 906.552
R369 C:F138 C:F70 251.979
R37 net020:F85 net020:F29 469.356
R370 C:F138 C:F66 71.7144
R371 C:F158 C:F142 15339.6
R372 C:F158 C:F86 81.544
R373 C:F158 C:F74 4255.03
R374 C:F158 C:F70 14609.1
R375 C:F158 C:F66 20888.7
R376 C:F142 C:F86 9686.93
R377 C:F142 C:F74 324.743
R378 C:F142 C:F70 90.2633
R379 C:F142 C:F66 251.979
R38 net020:F85 net020:F21 483.084
R380 C:F74 C:F86 4660.27
R381 C:F74 C:F70 309.279
R382 C:F74 C:F66 863.383
R383 C:F86 C:F70 16000.5
R384 C:F66 C:F70 239.98
R385 gnd gnd 0.001
R386 gnd gnd 9.33555
R387 gnd gnd 11.0541
R388 gnd gnd 6.13363
R389 gnd gnd 0.001
R39 net020:F85 net020:F19 494.423
R390 gnd gnd 3312.73
R391 gnd gnd 3290.55
R392 gnd gnd 3306.56
R393 gnd gnd 3305.35
R394 gnd gnd 40.0392
R395 gnd gnd 40.0392
R396 gnd gnd 39.7711
R397 gnd gnd 39.9646
R398 gnd gnd 39.95
R399 gnd gnd 37.5465
R4 net020:F53 net020:F61 349.846
R40 net020:F19 net020:F51 385.218
R400 gnd gnd 0.001
R401 gnd gnd 3305.35
R402 gnd gnd 3283.22
R403 gnd gnd 3299.19
R404 gnd gnd 0.001
R405 gnd gnd 3306.56
R406 gnd gnd 3284.42
R407 gnd gnd 0.001
R408 gnd gnd 3290.55
R409 gnd gnd 0.001
R41 net020:F19 net020:F37 355.07
R410 gnd gnd 0.001
R42 net020:F19 net020:F29 322.282
R43 net020:F19 net020:F21 288.502
R44 net020:F21 net020:F51 376.383
R45 net020:F21 net020:F37 346.926
R46 net020:F21 net020:F29 330.841
R47 net020:F21 net020:F27 0.001
R48 net020:F29 net020:F51 365.688
R49 net020:F29 net020:F37 337.068
R5 net020:F53 net020:F59 0.001
R50 net020:F29 net020:F35 0.001
R51 net020:F37 net020:F51 347.778
R52 net020:F37 net020:F43 0.001
R53 net020:F51 net020:F45 0.001
R54 net0158:F135 net0158:F129 0.001
R55 net0158:F135 net0158:F127 211.954
R56 net0158:F135 net0158:F119 224.686
R57 net0158:F135 net0158:F111 235.085
R58 net0158:F135 net0158:F103 242.47
R59 net0158:F135 net0158:F95 246.309
R6 net020:F53 net020:F51 372.524
R60 net0158:F119 net0158:F127 221.184
R61 net0158:F119 net0158:F113 0.001
R62 net0158:F119 net0158:F111 224.374
R63 net0158:F119 net0158:F103 231.422
R64 net0158:F119 net0158:F95 235.085
R65 net0158:F95 net0158:F127 242.47
R66 net0158:F95 net0158:F111 224.686
R67 net0158:F95 net0158:F103 211.954
R68 net0158:F95 net0158:F89 0.001
R69 net0158:F103 net0158:F127 238.692
R7 net020:F53 net020:F37 377.957
R70 net0158:F103 net0158:F111 221.184
R71 net0158:F103 net0158:F97 0.001
R72 net0158:F111 net0158:F127 231.422
R73 net0158:F111 net0158:F105 0.001
R74 net0158:F127 net0158:F121 0.001
R75 Z Z:F6 0.001
R76 Z:F131 Z:F151 8144.79
R77 Z:F131 Z:F125 0.001
R78 Z:F131 Z:F123 1642.72
R79 Z:F131 Z:F109 1668.25
R8 net020:F53 net020:F29 397.42
R80 Z:F131 Z:F6 40.4724
R81 Z:F109 Z:F143 5626.3
R82 Z:F109 Z:F123 1023.03
R83 Z:F109 Z:F115 0.001
R84 Z:F109 Z:F6 42.4786
R85 Z:F143 Z:F137 0.001
R86 Z:F143 Z:F123 5540.17
R87 Z:F143 Z:F6 18.9132
R88 Z:F6 Z:F159 39.4547
R89 Z:F6 Z:F151 38.8507
R9 net020:F53 net020:F21 409.044
R90 Z:F6 Z:F123 41.8284
R91 Z:F6 Z:F81 40.6206
R92 Z:F6 Z:F73 39.9177
R93 Z:F6 Z:F65 38.8303
R94 Z:F151 Z:F159 2701.27
R95 Z:F151 Z:F145 0.001
R96 Z:F159 Z:F153 0.001
R97 Z:F123 Z:F117 0.001
R98 Z:F65 Z:F81 3353.55
R99 Z:F65 Z:F73 3295.52
.ENDS HS65_GS_OAI21X37


