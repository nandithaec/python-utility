

`timescale 1ns/100ps

module dff (q, d,clk);

input clk, d;
output q;
reg q;
always @(posedge clk) 
q = d;

endmodule

// Verilog
// c432
// Ninputs 36
// Noutputs 7
// NtotalGates 160
// NOT1 40
// NAND2 64
// NOR2 19
// AND9 3
// XOR2 18
// NAND4 14
// AND8 1
// NAND3 1

module c432 (PCN1,PCN4,PCN8,PCN11,PCN14,PCN17,PCN21,PCN24,PCN27,PCN30,
             PCN34,PCN37,PCN40,PCN43,PCN47,PCN50,PCN53,PCN56,PCN60,PCN63,
             PCN66,PCN69,PCN73,PCN76,PCN79,PCN82,PCN86,PCN89,PCN92,PCN95,
             PCN99,PCN102,PCN105,PCN108,PCN112,PCN115,PCN223,PCN329,PCN370,PCN421,PCN430,PCN431,PCN432);

input PCN1,PCN4,PCN8,PCN11,PCN14,PCN17,PCN21,PCN24,PCN27,PCN30,
      PCN34,PCN37,PCN40,PCN43,PCN47,PCN50,PCN53,PCN56,PCN60,PCN63,
      PCN66,PCN69,PCN73,PCN76,PCN79,PCN82,PCN86,PCN89,PCN92,PCN95,
      PCN99,PCN102,PCN105,PCN108,PCN112,PCN115;

output PCN223,PCN329,PCN370,PCN421,PCN430,PCN431,PCN432;

wire PCN118,PCN119,PCN122,PCN123,PCN126,PCN127,PCN130,PCN131,PCN134,PCN135,
     PCN138,PCN139,PCN142,PCN143,PCN146,PCN147,PCN150,PCN151,PCN154,PCN157,
     PCN158,PCN159,PCN162,PCN165,PCN168,PCN171,PCN174,PCN177,PCN180,PCN183,
     PCN184,PCN185,PCN186,PCN187,PCN188,PCN189,PCN190,PCN191,PCN192,PCN193,
     PCN194,PCN195,PCN196,PCN197,PCN198,PCN199,PCN203,PCN213,PCN224,PCN227,
     PCN230,PCN233,PCN236,PCN239,PCN242,PCN243,PCN246,PCN247,PCN250,PCN251,
     PCN254,PCN255,PCN256,PCN257,PCN258,PCN259,PCN260,PCN263,PCN264,PCN267,
     PCN270,PCN273,PCN276,PCN279,PCN282,PCN285,PCN288,PCN289,PCN290,PCN291,
     PCN292,PCN293,PCN294,PCN295,PCN296,PCN300,PCN301,PCN302,PCN303,PCN304,
     PCN305,PCN306,PCN307,PCN308,PCN309,PCN319,PCN330,PCN331,PCN332,PCN333,
     PCN334,PCN335,PCN336,PCN337,PCN338,PCN339,PCN340,PCN341,PCN342,PCN343,
     PCN344,PCN345,PCN346,PCN347,PCN348,PCN349,PCN350,PCN351,PCN352,PCN353,
     PCN354,PCN355,PCN356,PCN357,PCN360,PCN371,PCN372,PCN373,PCN374,PCN375,
     PCN376,PCN377,PCN378,PCN379,PCN380,PCN381,PCN386,PCN393,PCN399,PCN404,
     PCN407,PCN411,PCN414,PCN415,PCN416,PCN417,PCN418,PCN419,PCN420,PCN422,
     PCN425,PCN428,PCN429;

not NOT1_1 (PCN118, PCN1);
not NOT1_2 (PCN119, PCN4);
not NOT1_3 (PCN122, PCN11);
not NOT1_4 (PCN123, PCN17);
not NOT1_5 (PCN126, PCN24);
not NOT1_6 (PCN127, PCN30);
not NOT1_7 (PCN130, PCN37);
not NOT1_8 (PCN131, PCN43);
not NOT1_9 (PCN134, PCN50);
not NOT1_10 (PCN135, PCN56);
not NOT1_11 (PCN138, PCN63);
not NOT1_12 (PCN139, PCN69);
not NOT1_13 (PCN142, PCN76);
not NOT1_14 (PCN143, PCN82);
not NOT1_15 (PCN146, PCN89);
not NOT1_16 (PCN147, PCN95);
not NOT1_17 (PCN150, PCN102);
not NOT1_18 (PCN151, PCN108);
nand NAND2_19 (PCN154, PCN118, PCN4);
nor NOR2_20 (PCN157, PCN8, PCN119);
nor NOR2_21 (PCN158, PCN14, PCN119);
nand NAND2_22 (PCN159, PCN122, PCN17);
nand NAND2_23 (PCN162, PCN126, PCN30);
nand NAND2_24 (PCN165, PCN130, PCN43);
nand NAND2_25 (PCN168, PCN134, PCN56);
nand NAND2_26 (PCN171, PCN138, PCN69);
nand NAND2_27 (PCN174, PCN142, PCN82);
nand NAND2_28 (PCN177, PCN146, PCN95);
nand NAND2_29 (PCN180, PCN150, PCN108);
nor NOR2_30 (PCN183, PCN21, PCN123);
nor NOR2_31 (PCN184, PCN27, PCN123);
nor NOR2_32 (PCN185, PCN34, PCN127);
nor NOR2_33 (PCN186, PCN40, PCN127);
nor NOR2_34 (PCN187, PCN47, PCN131);
nor NOR2_35 (PCN188, PCN53, PCN131);
nor NOR2_36 (PCN189, PCN60, PCN135);
nor NOR2_37 (PCN190, PCN66, PCN135);
nor NOR2_38 (PCN191, PCN73, PCN139);
nor NOR2_39 (PCN192, PCN79, PCN139);
nor NOR2_40 (PCN193, PCN86, PCN143);
nor NOR2_41 (PCN194, PCN92, PCN143);
nor NOR2_42 (PCN195, PCN99, PCN147);
nor NOR2_43 (PCN196, PCN105, PCN147);
nor NOR2_44 (PCN197, PCN112, PCN151);
nor NOR2_45 (PCN198, PCN115, PCN151);
and AND9_46 (PCN199, PCN154, PCN159, PCN162, PCN165, PCN168, PCN171, PCN174, PCN177, PCN180);
not NOT1_47 (PCN203, PCN199);
not NOT1_48 (PCN213, PCN199);
not NOT1_49 (PCN223, PCN199);
xor XOR2_50 (PCN224, PCN203, PCN154);
xor XOR2_51 (PCN227, PCN203, PCN159);
xor XOR2_52 (PCN230, PCN203, PCN162);
xor XOR2_53 (PCN233, PCN203, PCN165);
xor XOR2_54 (PCN236, PCN203, PCN168);
xor XOR2_55 (PCN239, PCN203, PCN171);
nand NAND2_56 (PCN242, PCN1, PCN213);
xor XOR2_57 (PCN243, PCN203, PCN174);
nand NAND2_58 (PCN246, PCN213, PCN11);
xor XOR2_59 (PCN247, PCN203, PCN177);
nand NAND2_60 (PCN250, PCN213, PCN24);
xor XOR2_61 (PCN251, PCN203, PCN180);
nand NAND2_62 (PCN254, PCN213, PCN37);
nand NAND2_63 (PCN255, PCN213, PCN50);
nand NAND2_64 (PCN256, PCN213, PCN63);
nand NAND2_65 (PCN257, PCN213, PCN76);
nand NAND2_66 (PCN258, PCN213, PCN89);
nand NAND2_67 (PCN259, PCN213, PCN102);
nand NAND2_68 (PCN260, PCN224, PCN157);
nand NAND2_69 (PCN263, PCN224, PCN158);
nand NAND2_70 (PCN264, PCN227, PCN183);
nand NAND2_71 (PCN267, PCN230, PCN185);
nand NAND2_72 (PCN270, PCN233, PCN187);
nand NAND2_73 (PCN273, PCN236, PCN189);
nand NAND2_74 (PCN276, PCN239, PCN191);
nand NAND2_75 (PCN279, PCN243, PCN193);
nand NAND2_76 (PCN282, PCN247, PCN195);
nand NAND2_77 (PCN285, PCN251, PCN197);
nand NAND2_78 (PCN288, PCN227, PCN184);
nand NAND2_79 (PCN289, PCN230, PCN186);
nand NAND2_80 (PCN290, PCN233, PCN188);
nand NAND2_81 (PCN291, PCN236, PCN190);
nand NAND2_82 (PCN292, PCN239, PCN192);
nand NAND2_83 (PCN293, PCN243, PCN194);
nand NAND2_84 (PCN294, PCN247, PCN196);
nand NAND2_85 (PCN295, PCN251, PCN198);
and AND9_86 (PCN296, PCN260, PCN264, PCN267, PCN270, PCN273, PCN276, PCN279, PCN282, PCN285);
not NOT1_87 (PCN300, PCN263);
not NOT1_88 (PCN301, PCN288);
not NOT1_89 (PCN302, PCN289);
not NOT1_90 (PCN303, PCN290);
not NOT1_91 (PCN304, PCN291);
not NOT1_92 (PCN305, PCN292);
not NOT1_93 (PCN306, PCN293);
not NOT1_94 (PCN307, PCN294);
not NOT1_95 (PCN308, PCN295);
not NOT1_96 (PCN309, PCN296);
not NOT1_97 (PCN319, PCN296);
not NOT1_98 (PCN329, PCN296);
xor XOR2_99 (PCN330, PCN309, PCN260);
xor XOR2_100 (PCN331, PCN309, PCN264);
xor XOR2_101 (PCN332, PCN309, PCN267);
xor XOR2_102 (PCN333, PCN309, PCN270);
nand NAND2_103 (PCN334, PCN8, PCN319);
xor XOR2_104 (PCN335, PCN309, PCN273);
nand NAND2_105 (PCN336, PCN319, PCN21);
xor XOR2_106 (PCN337, PCN309, PCN276);
nand NAND2_107 (PCN338, PCN319, PCN34);
xor XOR2_108 (PCN339, PCN309, PCN279);
nand NAND2_109 (PCN340, PCN319, PCN47);
xor XOR2_110 (PCN341, PCN309, PCN282);
nand NAND2_111 (PCN342, PCN319, PCN60);
xor XOR2_112 (PCN343, PCN309, PCN285);
nand NAND2_113 (PCN344, PCN319, PCN73);
nand NAND2_114 (PCN345, PCN319, PCN86);
nand NAND2_115 (PCN346, PCN319, PCN99);
nand NAND2_116 (PCN347, PCN319, PCN112);
nand NAND2_117 (PCN348, PCN330, PCN300);
nand NAND2_118 (PCN349, PCN331, PCN301);
nand NAND2_119 (PCN350, PCN332, PCN302);
nand NAND2_120 (PCN351, PCN333, PCN303);
nand NAND2_121 (PCN352, PCN335, PCN304);
nand NAND2_122 (PCN353, PCN337, PCN305);
nand NAND2_123 (PCN354, PCN339, PCN306);
nand NAND2_124 (PCN355, PCN341, PCN307);
nand NAND2_125 (PCN356, PCN343, PCN308);
and AND9_126 (PCN357, PCN348, PCN349, PCN350, PCN351, PCN352, PCN353, PCN354, PCN355, PCN356);
not NOT1_127 (PCN360, PCN357);
not NOT1_128 (PCN370, PCN357);
nand NAND2_129 (PCN371, PCN14, PCN360);
nand NAND2_130 (PCN372, PCN360, PCN27);
nand NAND2_131 (PCN373, PCN360, PCN40);
nand NAND2_132 (PCN374, PCN360, PCN53);
nand NAND2_133 (PCN375, PCN360, PCN66);
nand NAND2_134 (PCN376, PCN360, PCN79);
nand NAND2_135 (PCN377, PCN360, PCN92);
nand NAND2_136 (PCN378, PCN360, PCN105);
nand NAND2_137 (PCN379, PCN360, PCN115);
nand NAND4_138 (PCN380, PCN4, PCN242, PCN334, PCN371);
nand NAND4_139 (PCN381, PCN246, PCN336, PCN372, PCN17);
nand NAND4_140 (PCN386, PCN250, PCN338, PCN373, PCN30);
nand NAND4_141 (PCN393, PCN254, PCN340, PCN374, PCN43);
nand NAND4_142 (PCN399, PCN255, PCN342, PCN375, PCN56);
nand NAND4_143 (PCN404, PCN256, PCN344, PCN376, PCN69);
nand NAND4_144 (PCN407, PCN257, PCN345, PCN377, PCN82);
nand NAND4_145 (PCN411, PCN258, PCN346, PCN378, PCN95);
nand NAND4_146 (PCN414, PCN259, PCN347, PCN379, PCN108);
not NOT1_147 (PCN415, PCN380);
and AND8_148 (PCN416, PCN381, PCN386, PCN393, PCN399, PCN404, PCN407, PCN411, PCN414);
not NOT1_149 (PCN417, PCN393);
not NOT1_150 (PCN418, PCN404);
not NOT1_151 (PCN419, PCN407);
not NOT1_152 (PCN420, PCN411);
nor NOR2_153 (PCN421, PCN415, PCN416);
nand NAND2_154 (PCN422, PCN386, PCN417);
nand NAND4_155 (PCN425, PCN386, PCN393, PCN418, PCN399);
nand NAND3_156 (PCN428, PCN399, PCN393, PCN419);
nand NAND4_157 (PCN429, PCN386, PCN393, PCN407, PCN420);
nand NAND4_158 (PCN430, PCN381, PCN386, PCN422, PCN399);
nand NAND4_159 (PCN431, PCN381, PCN386, PCN425, PCN428);
nand NAND4_160 (PCN432, PCN381, PCN422, PCN425, PCN429);


endmodule



module c432_clk_ipFF (clk,PCN1,PCN4,PCN8,PCN11,PCN14,PCN17,PCN21,PCN24,PCN27,PCN30,
             PCN34,PCN37,PCN40,PCN43,PCN47,PCN50,PCN53,PCN56,PCN60,PCN63,
             PCN66,PCN69,PCN73,PCN76,PCN79,PCN82,PCN86,PCN89,PCN92,PCN95,
             PCN99,PCN102,PCN105,PCN108,PCN112,PCN115,Qout_PCN_223,Qout_PCN_329,Qout_PCN_370,Qout_PCN_421,
             Qout_PCN_430,Qout_PCN_431,Qout_PCN_432);

input clk,PCN1,PCN4,PCN8,PCN11,PCN14,PCN17,PCN21,PCN24,PCN27,PCN30,
      PCN34,PCN37,PCN40,PCN43,PCN47,PCN50,PCN53,PCN56,PCN60,PCN63,
      PCN66,PCN69,PCN73,PCN76,PCN79,PCN82,PCN86,PCN89,PCN92,PCN95,
      PCN99,PCN102,PCN105,PCN108,PCN112,PCN115;

output Qout_PCN_223,Qout_PCN_329,Qout_PCN_370,Qout_PCN_421,Qout_PCN_430,Qout_PCN_431,Qout_PCN_432;

wire PCN118,PCN119,PCN122,PCN123,PCN126,PCN127,PCN130,PCN131,PCN134,PCN135,
     PCN138,PCN139,PCN142,PCN143,PCN146,PCN147,PCN150,PCN151,PCN154,PCN157,
     PCN158,PCN159,PCN162,PCN165,PCN168,PCN171,PCN174,PCN177,PCN180,PCN183,
     PCN184,PCN185,PCN186,PCN187,PCN188,PCN189,PCN190,PCN191,PCN192,PCN193,
     PCN194,PCN195,PCN196,PCN197,PCN198,PCN199,PCN203,PCN213,PCN224,PCN227,
     PCN230,PCN233,PCN236,PCN239,PCN242,PCN243,PCN246,PCN247,PCN250,PCN251,
     PCN254,PCN255,PCN256,PCN257,PCN258,PCN259,PCN260,PCN263,PCN264,PCN267,
     PCN270,PCN273,PCN276,PCN279,PCN282,PCN285,PCN288,PCN289,PCN290,PCN291,
     PCN292,PCN293,PCN294,PCN295,PCN296,PCN300,PCN301,PCN302,PCN303,PCN304,
     PCN305,PCN306,PCN307,PCN308,PCN309,PCN319,PCN330,PCN331,PCN332,PCN333,
     PCN334,PCN335,PCN336,PCN337,PCN338,PCN339,PCN340,PCN341,PCN342,PCN343,
     PCN344,PCN345,PCN346,PCN347,PCN348,PCN349,PCN350,PCN351,PCN352,PCN353,
     PCN354,PCN355,PCN356,PCN357,PCN360,PCN371,PCN372,PCN373,PCN374,PCN375,
     PCN376,PCN377,PCN378,PCN379,PCN380,PCN381,PCN386,PCN393,PCN399,PCN404,
     PCN407,PCN411,PCN414,PCN415,PCN416,PCN417,PCN418,PCN419,PCN420,PCN422,
     PCN425,PCN428,PCN429;




 c432 C_0(INP_PCN1,INP_PCN4,INP_PCN8,INP_PCN11,INP_PCN14,INP_PCN17,INP_PCN21,INP_PCN24,INP_PCN27,INP_PCN30,
             INP_PCN34,INP_PCN37,INP_PCN40,INP_PCN43,INP_PCN47,INP_PCN50,INP_PCN53,INP_PCN56,INP_PCN60,INP_PCN63,
             INP_PCN66,INP_PCN69,INP_PCN73,INP_PCN76,INP_PCN79,INP_PCN82,INP_PCN86,INP_PCN89,INP_PCN92,INP_PCN95,
             INP_PCN99,INP_PCN102,INP_PCN105,INP_PCN108,INP_PCN112,INP_PCN115,DPCN_223,DPCN_329,DPCN_370,DPCN_421,
             DPCN_430,DPCN_431,DPCN_432);
	
	
//Input FFs
dff iDFF_1( INP_PCN1, PCN1, clk);
dff iDFF_2( INP_PCN4, PCN4, clk);
dff iDFF_3( INP_PCN8, PCN8, clk);
dff iDFF_4( INP_PCN11,PCN11, clk);
dff iDFF_5( INP_PCN14,PCN14, clk);
dff iDFF_6( INP_PCN17,PCN17, clk);
dff iDFF_7( INP_PCN21,PCN21, clk);
dff iDFF_8( INP_PCN24,PCN24, clk);
dff iDFF_9( INP_PCN27,PCN27, clk);
dff iDFF_10(INP_PCN30,PCN30, clk);
dff iDFF_12(INP_PCN34, PCN34, clk);
dff iDFF_13(INP_PCN37, PCN37, clk);
dff iDFF_14(INP_PCN40, PCN40, clk);
dff iDFF_15(INP_PCN43, PCN43, clk);
dff iDFF_16(INP_PCN47, PCN47, clk);
dff iDFF_17(INP_PCN50, PCN50, clk);
dff iDFF_18(INP_PCN53, PCN53, clk);
dff iDFF_19(INP_PCN56, PCN56, clk);
dff iDFF_20(INP_PCN60, PCN60, clk);
dff iDFF_21(INP_PCN63, PCN63, clk);
dff iDFF_23(INP_PCN66, PCN66, clk);
dff iDFF_24(INP_PCN69, PCN69, clk);
dff iDFF_25(INP_PCN73, PCN73, clk);
dff iDFF_26(INP_PCN76, PCN76, clk);
dff iDFF_27(INP_PCN79, PCN79, clk);
dff iDFF_28(INP_PCN82, PCN82, clk);
dff iDFF_29(INP_PCN86, PCN86, clk);
dff iDFF_30(INP_PCN89, PCN89, clk);
dff iDFF_31(INP_PCN92, PCN92, clk);
dff iDFF_32(INP_PCN95, PCN95, clk);
dff iDFF_34(INP_PCN99, PCN99, clk);
dff iDFF_35(INP_PCN102,PCN102, clk); 
dff iDFF_36(INP_PCN105,PCN105, clk);
dff iDFF_37(INP_PCN108,PCN108, clk); 
dff iDFF_38(INP_PCN112,PCN112, clk); 
dff iDFF_39(INP_PCN115,PCN115, clk); 


//Intermediate FFs
dff DFF_1(Qout_PCN_223,DPCN_223,clk);
dff DFF_2(Qout_PCN_329,DPCN_329,clk);
dff DFF_3(Qout_PCN_370,DPCN_370,clk);
dff DFF_4(Qout_PCN_421,DPCN_421,clk);
dff DFF_5(Qout_PCN_430,DPCN_430,clk);
dff DFF_6(Qout_PCN_431,DPCN_431,clk);
dff DFF_7(Qout_PCN_432,DPCN_432,clk);



endmodule



