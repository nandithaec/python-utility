
`timescale 1ns/100ps

module dff (q, d,clk);

input clk, d;
output q;
reg q;
always @(posedge clk) 
q = d;

endmodule

//32 outputs, 41 inputs
module c1355 (PGG1,PGG10,PGG11,PGG12,PGG13,PGG1324,PGG1325,PGG1326,PGG1327,PGG1328,PGG1329,PGG1330,
  PGG1331,PGG1332,PGG1333,PGG1334,PGG1335,PGG1336,PGG1337,PGG1338,PGG1339,PGG1340,PGG1341,PGG1342,
  PGG1343,PGG1344,PGG1345,PGG1346,PGG1347,PGG1348,PGG1349,PGG1350,PGG1351,PGG1352,PGG1353,PGG1354,
  PGG1355,PGG14,PGG15,PGG16,PGG17,PGG18,PGG19,PGG2,PGG20,PGG21,PGG22,PGG23,PGG24,PGG25,PGG26,PGG27,PGG28,PGG29,PGG3,
  PGG30,PGG31,PGG32,PGG33,PGG34,PGG35,PGG36,PGG37,PGG38,PGG39,PGG4,PGG40,PGG41,PGG5,PGG6,PGG7,PGG8,PGG9);

input PGG1,PGG2,PGG3,PGG4,PGG5,PGG6,PGG7,PGG8,PGG9,PGG10,PGG11,PGG12,PGG13,PGG14,PGG15,PGG16,PGG17,PGG18,PGG19,PGG20,
  PGG21,PGG22,PGG23,PGG24,PGG25,PGG26,PGG27,PGG28,PGG29,PGG30,PGG31,PGG32,PGG33,PGG34,PGG35,PGG36,PGG37,PGG38,PGG39,
  PGG40,PGG41;

output PGG1324,PGG1325,PGG1326,PGG1327,PGG1328,PGG1329,PGG1330,PGG1331,PGG1332,PGG1333,PGG1334,PGG1335,
  PGG1336,PGG1337,PGG1338,PGG1339,PGG1340,PGG1341,PGG1342,PGG1343,PGG1344,PGG1345,PGG1346,PGG1347,
  PGG1348,PGG1349,PGG1350,PGG1351,PGG1352,PGG1353,PGG1354,PGG1355;

  wire PGG242,PGG245,PGG248,PGG251,PGG254,PGG257,PGG260,PGG263,PGG266,PGG269,PGG272,PGG275,PGG278,PGG281,
    PGG284,PGG287,PGG290,PGG293,PGG296,PGG299,PGG302,PGG305,PGG308,PGG311,PGG314,PGG317,PGG320,PGG323,PGG326,
    PGG329,PGG332,PGG335,PGG338,PGG341,PGG344,PGG347,PGG350,PGG353,PGG356,PGG359,PGG362,PGG363,PGG364,PGG365,
    PGG366,PGG367,PGG368,PGG369,PGG370,PGG371,PGG372,PGG373,PGG374,PGG375,PGG376,PGG377,PGG378,PGG379,PGG380,
    PGG381,PGG382,PGG383,PGG384,PGG385,PGG386,PGG387,PGG388,PGG389,PGG390,PGG391,PGG392,PGG393,PGG394,PGG395,
    PGG396,PGG397,PGG398,PGG399,PGG400,PGG401,PGG402,PGG403,PGG404,PGG405,PGG406,PGG407,PGG408,PGG409,PGG410,
    PGG411,PGG412,PGG413,PGG414,PGG415,PGG416,PGG417,PGG418,PGG419,PGG420,PGG421,PGG422,PGG423,PGG424,PGG425,
    PGG426,PGG429,PGG432,PGG435,PGG438,PGG441,PGG444,PGG447,PGG450,PGG453,PGG456,PGG459,PGG462,PGG465,PGG468,
    PGG471,PGG474,PGG477,PGG480,PGG483,PGG486,PGG489,PGG492,PGG495,PGG498,PGG501,PGG504,PGG507,PGG510,PGG513,
    PGG516,PGG519,PGG522,PGG525,PGG528,PGG531,PGG534,PGG537,PGG540,PGG543,PGG546,PGG549,PGG552,PGG555,PGG558,
    PGG561,PGG564,PGG567,PGG570,PGG571,PGG572,PGG573,PGG574,PGG575,PGG576,PGG577,PGG578,PGG579,PGG580,PGG581,
    PGG582,PGG583,PGG584,PGG585,PGG586,PGG587,PGG588,PGG589,PGG590,PGG591,PGG592,PGG593,PGG594,PGG595,PGG596,
    PGG597,PGG598,PGG599,PGG600,PGG601,PGG602,PGG607,PGG612,PGG617,PGG622,PGG627,PGG632,PGG637,PGG642,PGG645,
    PGG648,PGG651,PGG654,PGG657,PGG660,PGG663,PGG666,PGG669,PGG672,PGG675,PGG678,PGG681,PGG684,PGG687,PGG690,
    PGG691,PGG692,PGG693,PGG694,PGG695,PGG696,PGG697,PGG698,PGG699,PGG700,PGG701,PGG702,PGG703,PGG704,PGG705,
    PGG706,PGG709,PGG712,PGG715,PGG718,PGG721,PGG724,PGG727,PGG730,PGG733,PGG736,PGG739,PGG742,PGG745,PGG748,
    PGG751,PGG754,PGG755,PGG756,PGG757,PGG758,PGG759,PGG760,PGG761,PGG762,PGG763,PGG764,PGG765,PGG766,PGG767,
    PGG768,PGG769,PGG770,PGG773,PGG776,PGG779,PGG782,PGG785,PGG788,PGG791,PGG794,PGG797,PGG800,PGG803,PGG806,
    PGG809,PGG812,PGG815,PGG818,PGG819,PGG820,PGG821,PGG822,PGG823,PGG824,PGG825,PGG826,PGG827,PGG828,PGG829,
    PGG830,PGG831,PGG832,PGG833,PGG834,PGG847,PGG860,PGG873,PGG886,PGG899,PGG912,PGG925,PGG938,PGG939,PGG940,
    PGG941,PGG942,PGG943,PGG944,PGG945,PGG946,PGG947,PGG948,PGG949,PGG950,PGG951,PGG952,PGG953,PGG954,PGG955,
    PGG956,PGG957,PGG958,PGG959,PGG960,PGG961,PGG962,PGG963,PGG964,PGG965,PGG966,PGG967,PGG968,PGG969,PGG970,
    PGG971,PGG972,PGG973,PGG974,PGG975,PGG976,PGG977,PGG978,PGG979,PGG980,PGG981,PGG982,PGG983,PGG984,PGG985,
    PGG986,PGG991,PGG996,PGG1001,PGG1006,PGG1011,PGG1016,PGG1021,PGG1026,PGG1031,PGG1036,PGG1039,PGG1042,
    PGG1045,PGG1048,PGG1051,PGG1054,PGG1057,PGG1060,PGG1063,PGG1066,PGG1069,PGG1072,PGG1075,PGG1078,
    PGG1081,PGG1084,PGG1087,PGG1090,PGG1093,PGG1096,PGG1099,PGG1102,PGG1105,PGG1108,PGG1111,PGG1114,
    PGG1117,PGG1120,PGG1123,PGG1126,PGG1129,PGG1132,PGG1135,PGG1138,PGG1141,PGG1144,PGG1147,PGG1150,
    PGG1153,PGG1156,PGG1159,PGG1162,PGG1165,PGG1168,PGG1171,PGG1174,PGG1177,PGG1180,PGG1183,PGG1186,
    PGG1189,PGG1192,PGG1195,PGG1198,PGG1201,PGG1204,PGG1207,PGG1210,PGG1213,PGG1216,PGG1219,PGG1222,
    PGG1225,PGG1228,PGG1229,PGG1230,PGG1231,PGG1232,PGG1233,PGG1234,PGG1235,PGG1236,PGG1237,PGG1238,
    PGG1239,PGG1240,PGG1241,PGG1242,PGG1243,PGG1244,PGG1245,PGG1246,PGG1247,PGG1248,PGG1249,PGG1250,
    PGG1251,PGG1252,PGG1253,PGG1254,PGG1255,PGG1256,PGG1257,PGG1258,PGG1259,PGG1260,PGG1261,PGG1262,
    PGG1263,PGG1264,PGG1265,PGG1266,PGG1267,PGG1268,PGG1269,PGG1270,PGG1271,PGG1272,PGG1273,PGG1274,
    PGG1275,PGG1276,PGG1277,PGG1278,PGG1279,PGG1280,PGG1281,PGG1282,PGG1283,PGG1284,PGG1285,PGG1286,
    PGG1287,PGG1288,PGG1289,PGG1290,PGG1291,PGG1292,PGG1293,PGG1294,PGG1295,PGG1296,PGG1297,PGG1298,
    PGG1299,PGG1300,PGG1301,PGG1302,PGG1303,PGG1304,PGG1305,PGG1306,PGG1307,PGG1308,PGG1309,PGG1310,
    PGG1311,PGG1312,PGG1313,PGG1314,PGG1315,PGG1316,PGG1317,PGG1318,PGG1319,PGG1320,PGG1321,PGG1322,
    PGG1323;

  and AND2_0(PGG242,PGG33,PGG41);
  and AND2_1(PGG245,PGG34,PGG41);
  and AND2_2(PGG248,PGG35,PGG41);
  and AND2_3(PGG251,PGG36,PGG41);
  and AND2_4(PGG254,PGG37,PGG41);
  and AND2_5(PGG257,PGG38,PGG41);
  and AND2_6(PGG260,PGG39,PGG41);
  and AND2_7(PGG263,PGG40,PGG41);
  nand NAND2_0(PGG266,PGG1,PGG2);
  nand NAND2_1(PGG269,PGG3,PGG4);
  nand NAND2_2(PGG272,PGG5,PGG6);
  nand NAND2_3(PGG275,PGG7,PGG8);
  nand NAND2_4(PGG278,PGG9,PGG10);
  nand NAND2_5(PGG281,PGG11,PGG12);
  nand NAND2_6(PGG284,PGG13,PGG14);
  nand NAND2_7(PGG287,PGG15,PGG16);
  nand NAND2_8(PGG290,PGG17,PGG18);
  nand NAND2_9(PGG293,PGG19,PGG20);
  nand NAND2_10(PGG296,PGG21,PGG22);
  nand NAND2_11(PGG299,PGG23,PGG24);
  nand NAND2_12(PGG302,PGG25,PGG26);
  nand NAND2_13(PGG305,PGG27,PGG28);
  nand NAND2_14(PGG308,PGG29,PGG30);
  nand NAND2_15(PGG311,PGG31,PGG32);
  nand NAND2_16(PGG314,PGG1,PGG5);
  nand NAND2_17(PGG317,PGG9,PGG13);
  nand NAND2_18(PGG320,PGG2,PGG6);
  nand NAND2_19(PGG323,PGG10,PGG14);
  nand NAND2_20(PGG326,PGG3,PGG7);
  nand NAND2_21(PGG329,PGG11,PGG15);
  nand NAND2_22(PGG332,PGG4,PGG8);
  nand NAND2_23(PGG335,PGG12,PGG16);
  nand NAND2_24(PGG338,PGG17,PGG21);
  nand NAND2_25(PGG341,PGG25,PGG29);
  nand NAND2_26(PGG344,PGG18,PGG22);
  nand NAND2_27(PGG347,PGG26,PGG30);
  nand NAND2_28(PGG350,PGG19,PGG23);
  nand NAND2_29(PGG353,PGG27,PGG31);
  nand NAND2_30(PGG356,PGG20,PGG24);
  nand NAND2_31(PGG359,PGG28,PGG32);
  nand NAND2_32(PGG362,PGG1,PGG266);
  nand NAND2_33(PGG363,PGG2,PGG266);
  nand NAND2_34(PGG364,PGG3,PGG269);
  nand NAND2_35(PGG365,PGG4,PGG269);
  nand NAND2_36(PGG366,PGG5,PGG272);
  nand NAND2_37(PGG367,PGG6,PGG272);
  nand NAND2_38(PGG368,PGG7,PGG275);
  nand NAND2_39(PGG369,PGG8,PGG275);
  nand NAND2_40(PGG370,PGG9,PGG278);
  nand NAND2_41(PGG371,PGG10,PGG278);
  nand NAND2_42(PGG372,PGG11,PGG281);
  nand NAND2_43(PGG373,PGG12,PGG281);
  nand NAND2_44(PGG374,PGG13,PGG284);
  nand NAND2_45(PGG375,PGG14,PGG284);
  nand NAND2_46(PGG376,PGG15,PGG287);
  nand NAND2_47(PGG377,PGG16,PGG287);
  nand NAND2_48(PGG378,PGG17,PGG290);
  nand NAND2_49(PGG379,PGG18,PGG290);
  nand NAND2_50(PGG380,PGG19,PGG293);
  nand NAND2_51(PGG381,PGG20,PGG293);
  nand NAND2_52(PGG382,PGG21,PGG296);
  nand NAND2_53(PGG383,PGG22,PGG296);
  nand NAND2_54(PGG384,PGG23,PGG299);
  nand NAND2_55(PGG385,PGG24,PGG299);
  nand NAND2_56(PGG386,PGG25,PGG302);
  nand NAND2_57(PGG387,PGG26,PGG302);
  nand NAND2_58(PGG388,PGG27,PGG305);
  nand NAND2_59(PGG389,PGG28,PGG305);
  nand NAND2_60(PGG390,PGG29,PGG308);
  nand NAND2_61(PGG391,PGG30,PGG308);
  nand NAND2_62(PGG392,PGG31,PGG311);
  nand NAND2_63(PGG393,PGG32,PGG311);
  nand NAND2_64(PGG394,PGG1,PGG314);
  nand NAND2_65(PGG395,PGG5,PGG314);
  nand NAND2_66(PGG396,PGG9,PGG317);
  nand NAND2_67(PGG397,PGG13,PGG317);
  nand NAND2_68(PGG398,PGG2,PGG320);
  nand NAND2_69(PGG399,PGG6,PGG320);
  nand NAND2_70(PGG400,PGG10,PGG323);
  nand NAND2_71(PGG401,PGG14,PGG323);
  nand NAND2_72(PGG402,PGG3,PGG326);
  nand NAND2_73(PGG403,PGG7,PGG326);
  nand NAND2_74(PGG404,PGG11,PGG329);
  nand NAND2_75(PGG405,PGG15,PGG329);
  nand NAND2_76(PGG406,PGG4,PGG332);
  nand NAND2_77(PGG407,PGG8,PGG332);
  nand NAND2_78(PGG408,PGG12,PGG335);
  nand NAND2_79(PGG409,PGG16,PGG335);
  nand NAND2_80(PGG410,PGG17,PGG338);
  nand NAND2_81(PGG411,PGG21,PGG338);
  nand NAND2_82(PGG412,PGG25,PGG341);
  nand NAND2_83(PGG413,PGG29,PGG341);
  nand NAND2_84(PGG414,PGG18,PGG344);
  nand NAND2_85(PGG415,PGG22,PGG344);
  nand NAND2_86(PGG416,PGG26,PGG347);
  nand NAND2_87(PGG417,PGG30,PGG347);
  nand NAND2_88(PGG418,PGG19,PGG350);
  nand NAND2_89(PGG419,PGG23,PGG350);
  nand NAND2_90(PGG420,PGG27,PGG353);
  nand NAND2_91(PGG421,PGG31,PGG353);
  nand NAND2_92(PGG422,PGG20,PGG356);
  nand NAND2_93(PGG423,PGG24,PGG356);
  nand NAND2_94(PGG424,PGG28,PGG359);
  nand NAND2_95(PGG425,PGG32,PGG359);
  nand NAND2_96(PGG426,PGG362,PGG363);
  nand NAND2_97(PGG429,PGG364,PGG365);
  nand NAND2_98(PGG432,PGG366,PGG367);
  nand NAND2_99(PGG435,PGG368,PGG369);
  nand NAND2_100(PGG438,PGG370,PGG371);
  nand NAND2_101(PGG441,PGG372,PGG373);
  nand NAND2_102(PGG444,PGG374,PGG375);
  nand NAND2_103(PGG447,PGG376,PGG377);
  nand NAND2_104(PGG450,PGG378,PGG379);
  nand NAND2_105(PGG453,PGG380,PGG381);
  nand NAND2_106(PGG456,PGG382,PGG383);
  nand NAND2_107(PGG459,PGG384,PGG385);
  nand NAND2_108(PGG462,PGG386,PGG387);
  nand NAND2_109(PGG465,PGG388,PGG389);
  nand NAND2_110(PGG468,PGG390,PGG391);
  nand NAND2_111(PGG471,PGG392,PGG393);
  nand NAND2_112(PGG474,PGG394,PGG395);
  nand NAND2_113(PGG477,PGG396,PGG397);
  nand NAND2_114(PGG480,PGG398,PGG399);
  nand NAND2_115(PGG483,PGG400,PGG401);
  nand NAND2_116(PGG486,PGG402,PGG403);
  nand NAND2_117(PGG489,PGG404,PGG405);
  nand NAND2_118(PGG492,PGG406,PGG407);
  nand NAND2_119(PGG495,PGG408,PGG409);
  nand NAND2_120(PGG498,PGG410,PGG411);
  nand NAND2_121(PGG501,PGG412,PGG413);
  nand NAND2_122(PGG504,PGG414,PGG415);
  nand NAND2_123(PGG507,PGG416,PGG417);
  nand NAND2_124(PGG510,PGG418,PGG419);
  nand NAND2_125(PGG513,PGG420,PGG421);
  nand NAND2_126(PGG516,PGG422,PGG423);
  nand NAND2_127(PGG519,PGG424,PGG425);
  nand NAND2_128(PGG522,PGG426,PGG429);
  nand NAND2_129(PGG525,PGG432,PGG435);
  nand NAND2_130(PGG528,PGG438,PGG441);
  nand NAND2_131(PGG531,PGG444,PGG447);
  nand NAND2_132(PGG534,PGG450,PGG453);
  nand NAND2_133(PGG537,PGG456,PGG459);
  nand NAND2_134(PGG540,PGG462,PGG465);
  nand NAND2_135(PGG543,PGG468,PGG471);
  nand NAND2_136(PGG546,PGG474,PGG477);
  nand NAND2_137(PGG549,PGG480,PGG483);
  nand NAND2_138(PGG552,PGG486,PGG489);
  nand NAND2_139(PGG555,PGG492,PGG495);
  nand NAND2_140(PGG558,PGG498,PGG501);
  nand NAND2_141(PGG561,PGG504,PGG507);
  nand NAND2_142(PGG564,PGG510,PGG513);
  nand NAND2_143(PGG567,PGG516,PGG519);
  nand NAND2_144(PGG570,PGG426,PGG522);
  nand NAND2_145(PGG571,PGG429,PGG522);
  nand NAND2_146(PGG572,PGG432,PGG525);
  nand NAND2_147(PGG573,PGG435,PGG525);
  nand NAND2_148(PGG574,PGG438,PGG528);
  nand NAND2_149(PGG575,PGG441,PGG528);
  nand NAND2_150(PGG576,PGG444,PGG531);
  nand NAND2_151(PGG577,PGG447,PGG531);
  nand NAND2_152(PGG578,PGG450,PGG534);
  nand NAND2_153(PGG579,PGG453,PGG534);
  nand NAND2_154(PGG580,PGG456,PGG537);
  nand NAND2_155(PGG581,PGG459,PGG537);
  nand NAND2_156(PGG582,PGG462,PGG540);
  nand NAND2_157(PGG583,PGG465,PGG540);
  nand NAND2_158(PGG584,PGG468,PGG543);
  nand NAND2_159(PGG585,PGG471,PGG543);
  nand NAND2_160(PGG586,PGG474,PGG546);
  nand NAND2_161(PGG587,PGG477,PGG546);
  nand NAND2_162(PGG588,PGG480,PGG549);
  nand NAND2_163(PGG589,PGG483,PGG549);
  nand NAND2_164(PGG590,PGG486,PGG552);
  nand NAND2_165(PGG591,PGG489,PGG552);
  nand NAND2_166(PGG592,PGG492,PGG555);
  nand NAND2_167(PGG593,PGG495,PGG555);
  nand NAND2_168(PGG594,PGG498,PGG558);
  nand NAND2_169(PGG595,PGG501,PGG558);
  nand NAND2_170(PGG596,PGG504,PGG561);
  nand NAND2_171(PGG597,PGG507,PGG561);
  nand NAND2_172(PGG598,PGG510,PGG564);
  nand NAND2_173(PGG599,PGG513,PGG564);
  nand NAND2_174(PGG600,PGG516,PGG567);
  nand NAND2_175(PGG601,PGG519,PGG567);
  nand NAND2_176(PGG602,PGG570,PGG571);
  nand NAND2_177(PGG607,PGG572,PGG573);
  nand NAND2_178(PGG612,PGG574,PGG575);
  nand NAND2_179(PGG617,PGG576,PGG577);
  nand NAND2_180(PGG622,PGG578,PGG579);
  nand NAND2_181(PGG627,PGG580,PGG581);
  nand NAND2_182(PGG632,PGG582,PGG583);
  nand NAND2_183(PGG637,PGG584,PGG585);
  nand NAND2_184(PGG642,PGG586,PGG587);
  nand NAND2_185(PGG645,PGG588,PGG589);
  nand NAND2_186(PGG648,PGG590,PGG591);
  nand NAND2_187(PGG651,PGG592,PGG593);
  nand NAND2_188(PGG654,PGG594,PGG595);
  nand NAND2_189(PGG657,PGG596,PGG597);
  nand NAND2_190(PGG660,PGG598,PGG599);
  nand NAND2_191(PGG663,PGG600,PGG601);
  nand NAND2_192(PGG666,PGG602,PGG607);
  nand NAND2_193(PGG669,PGG612,PGG617);
  nand NAND2_194(PGG672,PGG602,PGG612);
  nand NAND2_195(PGG675,PGG607,PGG617);
  nand NAND2_196(PGG678,PGG622,PGG627);
  nand NAND2_197(PGG681,PGG632,PGG637);
  nand NAND2_198(PGG684,PGG622,PGG632);
  nand NAND2_199(PGG687,PGG627,PGG637);
  nand NAND2_200(PGG690,PGG602,PGG666);
  nand NAND2_201(PGG691,PGG607,PGG666);
  nand NAND2_202(PGG692,PGG612,PGG669);
  nand NAND2_203(PGG693,PGG617,PGG669);
  nand NAND2_204(PGG694,PGG602,PGG672);
  nand NAND2_205(PGG695,PGG612,PGG672);
  nand NAND2_206(PGG696,PGG607,PGG675);
  nand NAND2_207(PGG697,PGG617,PGG675);
  nand NAND2_208(PGG698,PGG622,PGG678);
  nand NAND2_209(PGG699,PGG627,PGG678);
  nand NAND2_210(PGG700,PGG632,PGG681);
  nand NAND2_211(PGG701,PGG637,PGG681);
  nand NAND2_212(PGG702,PGG622,PGG684);
  nand NAND2_213(PGG703,PGG632,PGG684);
  nand NAND2_214(PGG704,PGG627,PGG687);
  nand NAND2_215(PGG705,PGG637,PGG687);
  nand NAND2_216(PGG706,PGG690,PGG691);
  nand NAND2_217(PGG709,PGG692,PGG693);
  nand NAND2_218(PGG712,PGG694,PGG695);
  nand NAND2_219(PGG715,PGG696,PGG697);
  nand NAND2_220(PGG718,PGG698,PGG699);
  nand NAND2_221(PGG721,PGG700,PGG701);
  nand NAND2_222(PGG724,PGG702,PGG703);
  nand NAND2_223(PGG727,PGG704,PGG705);
  nand NAND2_224(PGG730,PGG242,PGG718);
  nand NAND2_225(PGG733,PGG245,PGG721);
  nand NAND2_226(PGG736,PGG248,PGG724);
  nand NAND2_227(PGG739,PGG251,PGG727);
  nand NAND2_228(PGG742,PGG254,PGG706);
  nand NAND2_229(PGG745,PGG257,PGG709);
  nand NAND2_230(PGG748,PGG260,PGG712);
  nand NAND2_231(PGG751,PGG263,PGG715);
  nand NAND2_232(PGG754,PGG242,PGG730);
  nand NAND2_233(PGG755,PGG718,PGG730);
  nand NAND2_234(PGG756,PGG245,PGG733);
  nand NAND2_235(PGG757,PGG721,PGG733);
  nand NAND2_236(PGG758,PGG248,PGG736);
  nand NAND2_237(PGG759,PGG724,PGG736);
  nand NAND2_238(PGG760,PGG251,PGG739);
  nand NAND2_239(PGG761,PGG727,PGG739);
  nand NAND2_240(PGG762,PGG254,PGG742);
  nand NAND2_241(PGG763,PGG706,PGG742);
  nand NAND2_242(PGG764,PGG257,PGG745);
  nand NAND2_243(PGG765,PGG709,PGG745);
  nand NAND2_244(PGG766,PGG260,PGG748);
  nand NAND2_245(PGG767,PGG712,PGG748);
  nand NAND2_246(PGG768,PGG263,PGG751);
  nand NAND2_247(PGG769,PGG715,PGG751);
  nand NAND2_248(PGG770,PGG754,PGG755);
  nand NAND2_249(PGG773,PGG756,PGG757);
  nand NAND2_250(PGG776,PGG758,PGG759);
  nand NAND2_251(PGG779,PGG760,PGG761);
  nand NAND2_252(PGG782,PGG762,PGG763);
  nand NAND2_253(PGG785,PGG764,PGG765);
  nand NAND2_254(PGG788,PGG766,PGG767);
  nand NAND2_255(PGG791,PGG768,PGG769);
  nand NAND2_256(PGG794,PGG642,PGG770);
  nand NAND2_257(PGG797,PGG645,PGG773);
  nand NAND2_258(PGG800,PGG648,PGG776);
  nand NAND2_259(PGG803,PGG651,PGG779);
  nand NAND2_260(PGG806,PGG654,PGG782);
  nand NAND2_261(PGG809,PGG657,PGG785);
  nand NAND2_262(PGG812,PGG660,PGG788);
  nand NAND2_263(PGG815,PGG663,PGG791);
  nand NAND2_264(PGG818,PGG642,PGG794);
  nand NAND2_265(PGG819,PGG770,PGG794);
  nand NAND2_266(PGG820,PGG645,PGG797);
  nand NAND2_267(PGG821,PGG773,PGG797);
  nand NAND2_268(PGG822,PGG648,PGG800);
  nand NAND2_269(PGG823,PGG776,PGG800);
  nand NAND2_270(PGG824,PGG651,PGG803);
  nand NAND2_271(PGG825,PGG779,PGG803);
  nand NAND2_272(PGG826,PGG654,PGG806);
  nand NAND2_273(PGG827,PGG782,PGG806);
  nand NAND2_274(PGG828,PGG657,PGG809);
  nand NAND2_275(PGG829,PGG785,PGG809);
  nand NAND2_276(PGG830,PGG660,PGG812);
  nand NAND2_277(PGG831,PGG788,PGG812);
  nand NAND2_278(PGG832,PGG663,PGG815);
  nand NAND2_279(PGG833,PGG791,PGG815);
  nand NAND2_280(PGG834,PGG818,PGG819);
  nand NAND2_281(PGG847,PGG820,PGG821);
  nand NAND2_282(PGG860,PGG822,PGG823);
  nand NAND2_283(PGG873,PGG824,PGG825);
  nand NAND2_284(PGG886,PGG828,PGG829);
  nand NAND2_285(PGG899,PGG832,PGG833);
  nand NAND2_286(PGG912,PGG830,PGG831);
  nand NAND2_287(PGG925,PGG826,PGG827);
  not NOT_0(PGG938,PGG834);
  not NOT_1(PGG939,PGG847);
  not NOT_2(PGG940,PGG860);
  not NOT_3(PGG941,PGG834);
  not NOT_4(PGG942,PGG847);
  not NOT_5(PGG943,PGG873);
  not NOT_6(PGG944,PGG834);
  not NOT_7(PGG945,PGG860);
  not NOT_8(PGG946,PGG873);
  not NOT_9(PGG947,PGG847);
  not NOT_10(PGG948,PGG860);
  not NOT_11(PGG949,PGG873);
  not NOT_12(PGG950,PGG886);
  not NOT_13(PGG951,PGG899);
  not NOT_14(PGG952,PGG886);
  not NOT_15(PGG953,PGG912);
  not NOT_16(PGG954,PGG925);
  not NOT_17(PGG955,PGG899);
  not NOT_18(PGG956,PGG925);
  not NOT_19(PGG957,PGG912);
  not NOT_20(PGG958,PGG925);
  not NOT_21(PGG959,PGG886);
  not NOT_22(PGG960,PGG912);
  not NOT_23(PGG961,PGG925);
  not NOT_24(PGG962,PGG886);
  not NOT_25(PGG963,PGG899);
  not NOT_26(PGG964,PGG925);
  not NOT_27(PGG965,PGG912);
  not NOT_28(PGG966,PGG899);
  not NOT_29(PGG967,PGG886);
  not NOT_30(PGG968,PGG912);
  not NOT_31(PGG969,PGG899);
  not NOT_32(PGG970,PGG847);
  not NOT_33(PGG971,PGG873);
  not NOT_34(PGG972,PGG847);
  not NOT_35(PGG973,PGG860);
  not NOT_36(PGG974,PGG834);
  not NOT_37(PGG975,PGG873);
  not NOT_38(PGG976,PGG834);
  not NOT_39(PGG977,PGG860);
  and AND4_0(PGG978,PGG938,PGG939,PGG940,PGG873);
  and AND4_1(PGG979,PGG941,PGG942,PGG860,PGG943);
  and AND4_2(PGG980,PGG944,PGG847,PGG945,PGG946);
  and AND4_3(PGG981,PGG834,PGG947,PGG948,PGG949);
  and AND4_4(PGG982,PGG958,PGG959,PGG960,PGG899);
  and AND4_5(PGG983,PGG961,PGG962,PGG912,PGG963);
  and AND4_6(PGG984,PGG964,PGG886,PGG965,PGG966);
  and AND4_7(PGG985,PGG925,PGG967,PGG968,PGG969);
  or OR4_0(PGG986,PGG978,PGG979,PGG980,PGG981);
  or OR4_1(PGG991,PGG982,PGG983,PGG984,PGG985);
  and AND5_0(PGG996,PGG925,PGG950,PGG912,PGG951,PGG986);
  and AND5_1(PGG1001,PGG925,PGG952,PGG953,PGG899,PGG986);
  and AND5_2(PGG1006,PGG954,PGG886,PGG912,PGG955,PGG986);
  and AND5_3(PGG1011,PGG956,PGG886,PGG957,PGG899,PGG986);
  and AND5_4(PGG1016,PGG834,PGG970,PGG860,PGG971,PGG991);
  and AND5_5(PGG1021,PGG834,PGG972,PGG973,PGG873,PGG991);
  and AND5_6(PGG1026,PGG974,PGG847,PGG860,PGG975,PGG991);
  and AND5_7(PGG1031,PGG976,PGG847,PGG977,PGG873,PGG991);
  and AND2_8(PGG1036,PGG834,PGG996);
  and AND2_9(PGG1039,PGG847,PGG996);
  and AND2_10(PGG1042,PGG860,PGG996);
  and AND2_11(PGG1045,PGG873,PGG996);
  and AND2_12(PGG1048,PGG834,PGG1001);
  and AND2_13(PGG1051,PGG847,PGG1001);
  and AND2_14(PGG1054,PGG860,PGG1001);
  and AND2_15(PGG1057,PGG873,PGG1001);
  and AND2_16(PGG1060,PGG834,PGG1006);
  and AND2_17(PGG1063,PGG847,PGG1006);
  and AND2_18(PGG1066,PGG860,PGG1006);
  and AND2_19(PGG1069,PGG873,PGG1006);
  and AND2_20(PGG1072,PGG834,PGG1011);
  and AND2_21(PGG1075,PGG847,PGG1011);
  and AND2_22(PGG1078,PGG860,PGG1011);
  and AND2_23(PGG1081,PGG873,PGG1011);
  and AND2_24(PGG1084,PGG925,PGG1016);
  and AND2_25(PGG1087,PGG886,PGG1016);
  and AND2_26(PGG1090,PGG912,PGG1016);
  and AND2_27(PGG1093,PGG899,PGG1016);
  and AND2_28(PGG1096,PGG925,PGG1021);
  and AND2_29(PGG1099,PGG886,PGG1021);
  and AND2_30(PGG1102,PGG912,PGG1021);
  and AND2_31(PGG1105,PGG899,PGG1021);
  and AND2_32(PGG1108,PGG925,PGG1026);
  and AND2_33(PGG1111,PGG886,PGG1026);
  and AND2_34(PGG1114,PGG912,PGG1026);
  and AND2_35(PGG1117,PGG899,PGG1026);
  and AND2_36(PGG1120,PGG925,PGG1031);
  and AND2_37(PGG1123,PGG886,PGG1031);
  and AND2_38(PGG1126,PGG912,PGG1031);
  and AND2_39(PGG1129,PGG899,PGG1031);
  nand NAND2_288(PGG1132,PGG1,PGG1036);
  nand NAND2_289(PGG1135,PGG2,PGG1039);
  nand NAND2_290(PGG1138,PGG3,PGG1042);
  nand NAND2_291(PGG1141,PGG4,PGG1045);
  nand NAND2_292(PGG1144,PGG5,PGG1048);
  nand NAND2_293(PGG1147,PGG6,PGG1051);
  nand NAND2_294(PGG1150,PGG7,PGG1054);
  nand NAND2_295(PGG1153,PGG8,PGG1057);
  nand NAND2_296(PGG1156,PGG9,PGG1060);
  nand NAND2_297(PGG1159,PGG10,PGG1063);
  nand NAND2_298(PGG1162,PGG11,PGG1066);
  nand NAND2_299(PGG1165,PGG12,PGG1069);
  nand NAND2_300(PGG1168,PGG13,PGG1072);
  nand NAND2_301(PGG1171,PGG14,PGG1075);
  nand NAND2_302(PGG1174,PGG15,PGG1078);
  nand NAND2_303(PGG1177,PGG16,PGG1081);
  nand NAND2_304(PGG1180,PGG17,PGG1084);
  nand NAND2_305(PGG1183,PGG18,PGG1087);
  nand NAND2_306(PGG1186,PGG19,PGG1090);
  nand NAND2_307(PGG1189,PGG20,PGG1093);
  nand NAND2_308(PGG1192,PGG21,PGG1096);
  nand NAND2_309(PGG1195,PGG22,PGG1099);
  nand NAND2_310(PGG1198,PGG23,PGG1102);
  nand NAND2_311(PGG1201,PGG24,PGG1105);
  nand NAND2_312(PGG1204,PGG25,PGG1108);
  nand NAND2_313(PGG1207,PGG26,PGG1111);
  nand NAND2_314(PGG1210,PGG27,PGG1114);
  nand NAND2_315(PGG1213,PGG28,PGG1117);
  nand NAND2_316(PGG1216,PGG29,PGG1120);
  nand NAND2_317(PGG1219,PGG30,PGG1123);
  nand NAND2_318(PGG1222,PGG31,PGG1126);
  nand NAND2_319(PGG1225,PGG32,PGG1129);
  nand NAND2_320(PGG1228,PGG1,PGG1132);
  nand NAND2_321(PGG1229,PGG1036,PGG1132);
  nand NAND2_322(PGG1230,PGG2,PGG1135);
  nand NAND2_323(PGG1231,PGG1039,PGG1135);
  nand NAND2_324(PGG1232,PGG3,PGG1138);
  nand NAND2_325(PGG1233,PGG1042,PGG1138);
  nand NAND2_326(PGG1234,PGG4,PGG1141);
  nand NAND2_327(PGG1235,PGG1045,PGG1141);
  nand NAND2_328(PGG1236,PGG5,PGG1144);
  nand NAND2_329(PGG1237,PGG1048,PGG1144);
  nand NAND2_330(PGG1238,PGG6,PGG1147);
  nand NAND2_331(PGG1239,PGG1051,PGG1147);
  nand NAND2_332(PGG1240,PGG7,PGG1150);
  nand NAND2_333(PGG1241,PGG1054,PGG1150);
  nand NAND2_334(PGG1242,PGG8,PGG1153);
  nand NAND2_335(PGG1243,PGG1057,PGG1153);
  nand NAND2_336(PGG1244,PGG9,PGG1156);
  nand NAND2_337(PGG1245,PGG1060,PGG1156);
  nand NAND2_338(PGG1246,PGG10,PGG1159);
  nand NAND2_339(PGG1247,PGG1063,PGG1159);
  nand NAND2_340(PGG1248,PGG11,PGG1162);
  nand NAND2_341(PGG1249,PGG1066,PGG1162);
  nand NAND2_342(PGG1250,PGG12,PGG1165);
  nand NAND2_343(PGG1251,PGG1069,PGG1165);
  nand NAND2_344(PGG1252,PGG13,PGG1168);
  nand NAND2_345(PGG1253,PGG1072,PGG1168);
  nand NAND2_346(PGG1254,PGG14,PGG1171);
  nand NAND2_347(PGG1255,PGG1075,PGG1171);
  nand NAND2_348(PGG1256,PGG15,PGG1174);
  nand NAND2_349(PGG1257,PGG1078,PGG1174);
  nand NAND2_350(PGG1258,PGG16,PGG1177);
  nand NAND2_351(PGG1259,PGG1081,PGG1177);
  nand NAND2_352(PGG1260,PGG17,PGG1180);
  nand NAND2_353(PGG1261,PGG1084,PGG1180);
  nand NAND2_354(PGG1262,PGG18,PGG1183);
  nand NAND2_355(PGG1263,PGG1087,PGG1183);
  nand NAND2_356(PGG1264,PGG19,PGG1186);
  nand NAND2_357(PGG1265,PGG1090,PGG1186);
  nand NAND2_358(PGG1266,PGG20,PGG1189);
  nand NAND2_359(PGG1267,PGG1093,PGG1189);
  nand NAND2_360(PGG1268,PGG21,PGG1192);
  nand NAND2_361(PGG1269,PGG1096,PGG1192);
  nand NAND2_362(PGG1270,PGG22,PGG1195);
  nand NAND2_363(PGG1271,PGG1099,PGG1195);
  nand NAND2_364(PGG1272,PGG23,PGG1198);
  nand NAND2_365(PGG1273,PGG1102,PGG1198);
  nand NAND2_366(PGG1274,PGG24,PGG1201);
  nand NAND2_367(PGG1275,PGG1105,PGG1201);
  nand NAND2_368(PGG1276,PGG25,PGG1204);
  nand NAND2_369(PGG1277,PGG1108,PGG1204);
  nand NAND2_370(PGG1278,PGG26,PGG1207);
  nand NAND2_371(PGG1279,PGG1111,PGG1207);
  nand NAND2_372(PGG1280,PGG27,PGG1210);
  nand NAND2_373(PGG1281,PGG1114,PGG1210);
  nand NAND2_374(PGG1282,PGG28,PGG1213);
  nand NAND2_375(PGG1283,PGG1117,PGG1213);
  nand NAND2_376(PGG1284,PGG29,PGG1216);
  nand NAND2_377(PGG1285,PGG1120,PGG1216);
  nand NAND2_378(PGG1286,PGG30,PGG1219);
  nand NAND2_379(PGG1287,PGG1123,PGG1219);
  nand NAND2_380(PGG1288,PGG31,PGG1222);
  nand NAND2_381(PGG1289,PGG1126,PGG1222);
  nand NAND2_382(PGG1290,PGG32,PGG1225);
  nand NAND2_383(PGG1291,PGG1129,PGG1225);
  nand NAND2_384(PGG1292,PGG1228,PGG1229);
  nand NAND2_385(PGG1293,PGG1230,PGG1231);
  nand NAND2_386(PGG1294,PGG1232,PGG1233);
  nand NAND2_387(PGG1295,PGG1234,PGG1235);
  nand NAND2_388(PGG1296,PGG1236,PGG1237);
  nand NAND2_389(PGG1297,PGG1238,PGG1239);
  nand NAND2_390(PGG1298,PGG1240,PGG1241);
  nand NAND2_391(PGG1299,PGG1242,PGG1243);
  nand NAND2_392(PGG1300,PGG1244,PGG1245);
  nand NAND2_393(PGG1301,PGG1246,PGG1247);
  nand NAND2_394(PGG1302,PGG1248,PGG1249);
  nand NAND2_395(PGG1303,PGG1250,PGG1251);
  nand NAND2_396(PGG1304,PGG1252,PGG1253);
  nand NAND2_397(PGG1305,PGG1254,PGG1255);
  nand NAND2_398(PGG1306,PGG1256,PGG1257);
  nand NAND2_399(PGG1307,PGG1258,PGG1259);
  nand NAND2_400(PGG1308,PGG1260,PGG1261);
  nand NAND2_401(PGG1309,PGG1262,PGG1263);
  nand NAND2_402(PGG1310,PGG1264,PGG1265);
  nand NAND2_403(PGG1311,PGG1266,PGG1267);
  nand NAND2_404(PGG1312,PGG1268,PGG1269);
  nand NAND2_405(PGG1313,PGG1270,PGG1271);
  nand NAND2_406(PGG1314,PGG1272,PGG1273);
  nand NAND2_407(PGG1315,PGG1274,PGG1275);
  nand NAND2_408(PGG1316,PGG1276,PGG1277);
  nand NAND2_409(PGG1317,PGG1278,PGG1279);
  nand NAND2_410(PGG1318,PGG1280,PGG1281);
  nand NAND2_411(PGG1319,PGG1282,PGG1283);
  nand NAND2_412(PGG1320,PGG1284,PGG1285);
  nand NAND2_413(PGG1321,PGG1286,PGG1287);
  nand NAND2_414(PGG1322,PGG1288,PGG1289);
  nand NAND2_415(PGG1323,PGG1290,PGG1291);
  not NOT_40(PGG1324,PGG1292);
  not NOT_41(PGG1325,PGG1293);
  not NOT_42(PGG1326,PGG1294);
  not NOT_43(PGG1327,PGG1295);
  not NOT_44(PGG1328,PGG1296);
  not NOT_45(PGG1329,PGG1297);
  not NOT_46(PGG1330,PGG1298);
  not NOT_47(PGG1331,PGG1299);
  not NOT_48(PGG1332,PGG1300);
  not NOT_49(PGG1333,PGG1301);
  not NOT_50(PGG1334,PGG1302);
  not NOT_51(PGG1335,PGG1303);
  not NOT_52(PGG1336,PGG1304);
  not NOT_53(PGG1337,PGG1305);
  not NOT_54(PGG1338,PGG1306);
  not NOT_55(PGG1339,PGG1307);
  not NOT_56(PGG1340,PGG1308);
  not NOT_57(PGG1341,PGG1309);
  not NOT_58(PGG1342,PGG1310);
  not NOT_59(PGG1343,PGG1311);
  not NOT_60(PGG1344,PGG1312);
  not NOT_61(PGG1345,PGG1313);
  not NOT_62(PGG1346,PGG1314);
  not NOT_63(PGG1347,PGG1315);
  not NOT_64(PGG1348,PGG1316);
  not NOT_65(PGG1349,PGG1317);
  not NOT_66(PGG1350,PGG1318);
  not NOT_67(PGG1351,PGG1319);
  not NOT_68(PGG1352,PGG1320);
  not NOT_69(PGG1353,PGG1321);
  not NOT_70(PGG1354,PGG1322);
  not NOT_71(PGG1355,PGG1323);

endmodule


module c1355_clk_ipFF (clk,PGG1,PGG10,PGG11,PGG12,PGG13,
	Q_PGG1324,Q_PGG1325,Q_PGG1326,Q_PGG1327,Q_PGG1328,Q_PGG1329,Q_PGG1330,
  Q_PGG1331,Q_PGG1332,Q_PGG1333,Q_PGG1334,Q_PGG1335,Q_PGG1336,Q_PGG1337,Q_PGG1338,Q_PGG1339,Q_PGG1340,Q_PGG1341,Q_PGG1342,
  Q_PGG1343,Q_PGG1344,Q_PGG1345,Q_PGG1346,Q_PGG1347,Q_PGG1348,Q_PGG1349,Q_PGG1350,Q_PGG1351,Q_PGG1352,Q_PGG1353,Q_PGG1354,
  Q_PGG1355,
	PGG14,PGG15,PGG16,PGG17,PGG18,PGG19,PGG2,PGG20,PGG21,PGG22,PGG23,PGG24,PGG25,PGG26,PGG27,PGG28,PGG29,PGG3,
  PGG30,PGG31,PGG32,PGG33,PGG34,PGG35,PGG36,PGG37,PGG38,PGG39,PGG4,PGG40,PGG41,PGG5,PGG6,PGG7,PGG8,PGG9);

input clk,PGG1,PGG2,PGG3,PGG4,PGG5,PGG6,PGG7,PGG8,PGG9,PGG10,PGG11,PGG12,PGG13,PGG14,PGG15,PGG16,PGG17,PGG18,PGG19,PGG20,
  PGG21,PGG22,PGG23,PGG24,PGG25,PGG26,PGG27,PGG28,PGG29,PGG30,PGG31,PGG32,PGG33,PGG34,PGG35,PGG36,PGG37,PGG38,PGG39,
  PGG40,PGG41;

output Q_PGG1324,Q_PGG1325,Q_PGG1326,Q_PGG1327,Q_PGG1328,Q_PGG1329,Q_PGG1330,
  Q_PGG1331,Q_PGG1332,Q_PGG1333,Q_PGG1334,Q_PGG1335,Q_PGG1336,Q_PGG1337,Q_PGG1338,Q_PGG1339,Q_PGG1340,Q_PGG1341,
  Q_PGG1342, Q_PGG1343,Q_PGG1344,Q_PGG1345,Q_PGG1346,Q_PGG1347,Q_PGG1348,Q_PGG1349,Q_PGG1350,Q_PGG1351,Q_PGG1352,
  Q_PGG1353, Q_PGG1354, Q_PGG1355;

c1355 c1 (INP_PGG1,INP_PGG10,INP_PGG11,INP_PGG12,INP_PGG13,PGG1324,PGG1325,PGG1326,PGG1327,PGG1328,PGG1329,PGG1330,
  PGG1331,PGG1332,PGG1333,PGG1334,PGG1335,PGG1336,PGG1337,PGG1338,PGG1339,PGG1340,PGG1341,PGG1342,
  PGG1343,PGG1344,PGG1345,PGG1346,PGG1347,PGG1348,PGG1349,PGG1350,PGG1351,PGG1352,PGG1353,PGG1354,
PGG1355,INP_PGG14,INP_PGG15,INP_PGG16,INP_PGG17,INP_PGG18,INP_PGG19,INP_PGG2,INP_PGG20,INP_PGG21,INP_PGG22,INP_PGG23,
  INP_PGG24,INP_PGG25,INP_PGG26,INP_PGG27,INP_PGG28,INP_PGG29,INP_PGG3,
  INP_PGG30,INP_PGG31,INP_PGG32,INP_PGG33,INP_PGG34,INP_PGG35,INP_PGG36,INP_PGG37,INP_PGG38,
  INP_PGG39,INP_PGG4,INP_PGG40,INP_PGG41,INP_PGG5,INP_PGG6,INP_PGG7,INP_PGG8,INP_PGG9);

//input FFs
dff iDFF_1(  INP_PGG1, PGG1, clk);
dff iDFF_2(  INP_PGG2, PGG2, clk);
dff iDFF_3(  INP_PGG3, PGG3, clk);
dff iDFF_4(  INP_PGG4, PGG4, clk);
dff iDFF_5(  INP_PGG5, PGG5, clk);
dff iDFF_6(  INP_PGG6, PGG6, clk);
dff iDFF_7(  INP_PGG7, PGG7, clk);
dff iDFF_8(  INP_PGG8, PGG8, clk);
dff iDFF_9(  INP_PGG9, PGG9, clk);
dff iDFF_10( INP_PGG10,PGG10, clk);
dff iDFF_11( INP_PGG11,PGG11, clk);
dff iDFF_12( INP_PGG12,PGG12, clk);
dff iDFF_13( INP_PGG13,PGG13, clk);
dff iDFF_14( INP_PGG14,PGG14, clk);
dff iDFF_15( INP_PGG15,PGG15, clk);
dff iDFF_16( INP_PGG16,PGG16, clk);
dff iDFF_17( INP_PGG17,PGG17, clk);
dff iDFF_18( INP_PGG18,PGG18, clk);
dff iDFF_19( INP_PGG19,PGG19, clk);
dff iDFF_20( INP_PGG20,PGG20, clk);
dff iDFF_21( INP_PGG21,PGG21, clk);
dff iDFF_22( INP_PGG22,PGG22, clk);
dff iDFF_23( INP_PGG23,PGG23, clk);
dff iDFF_24( INP_PGG24,PGG24, clk);
dff iDFF_25( INP_PGG25,PGG25, clk);
dff iDFF_26( INP_PGG26,PGG26, clk);
dff iDFF_27( INP_PGG27,PGG27, clk);
dff iDFF_28( INP_PGG28,PGG28, clk);
dff iDFF_29( INP_PGG29,PGG29, clk);
dff iDFF_30( INP_PGG30,PGG30, clk);
dff iDFF_31( INP_PGG31,PGG31, clk);
dff iDFF_32( INP_PGG32,PGG32, clk);
dff iDFF_33( INP_PGG33,PGG33, clk);
dff iDFF_34( INP_PGG34,PGG34, clk);
dff iDFF_35( INP_PGG35,PGG35, clk);
dff iDFF_36( INP_PGG36,PGG36, clk);
dff iDFF_37( INP_PGG37,PGG37, clk);
dff iDFF_38( INP_PGG38,PGG38, clk);
dff iDFF_39( INP_PGG39,PGG39, clk);
dff iDFF_40( INP_PGG40,PGG40, clk);
dff iDFF_41( INP_PGG41, PGG41, clk);


//output FFs
dff DFF_1   (Q_PGG1324, PGG1324,clk);
dff DFF_2   (Q_PGG1325, PGG1325,clk);
dff DFF_3   (Q_PGG1326, PGG1326,clk);
dff DFF_4   (Q_PGG1327, PGG1327,clk);
dff DFF_5   (Q_PGG1328, PGG1328,clk);
dff DFF_6   (Q_PGG1329, PGG1329,clk);
dff DFF_7   (Q_PGG1330, PGG1330,clk);
dff DFF_8   (Q_PGG1331, PGG1331,clk);
dff DFF_9   (Q_PGG1332, PGG1332,clk);
dff DFF_10   (Q_PGG1333, PGG1333,clk);
dff DFF_11   (Q_PGG1334, PGG1334,clk);
dff DFF_12   (Q_PGG1335, PGG1335,clk);
dff DFF_13   (Q_PGG1336, PGG1336,clk);
dff DFF_14   (Q_PGG1337, PGG1337,clk);
dff DFF_15   (Q_PGG1338, PGG1338,clk);
dff DFF_16   (Q_PGG1339, PGG1339,clk);
dff DFF_17   (Q_PGG1340, PGG1340,clk);
dff DFF_18   (Q_PGG1341, PGG1341,clk);
dff DFF_19   (Q_PGG1342, PGG1342,clk);
dff DFF_20   (Q_PGG1343, PGG1343,clk);
dff DFF_21   (Q_PGG1344, PGG1344,clk);
dff DFF_22   (Q_PGG1345, PGG1345,clk);
dff DFF_23   (Q_PGG1346, PGG1346,clk);
dff DFF_24   (Q_PGG1347, PGG1347,clk);
dff DFF_25   (Q_PGG1348, PGG1348,clk);
dff DFF_26   (Q_PGG1349, PGG1349,clk);
dff DFF_27   (Q_PGG1350, PGG1350,clk);
dff DFF_28   (Q_PGG1351, PGG1351,clk);
dff DFF_29   (Q_PGG1352, PGG1352,clk);
dff DFF_30   (Q_PGG1353, PGG1353,clk);
dff DFF_31   (Q_PGG1354, PGG1354,clk);
dff DFF_32   (Q_PGG1355, PGG1355,clk);


endmodule
