

`timescale 1ns/100ps

module dff (q, d,clk);

input clk, d;
output q;
reg q;
always @(posedge clk) 
q = d;

endmodule

// Verilog
// c1908
// Ninputs 33
// Noutputs 25
// NtotalGates 880
// NOT1 277
// NAND2 347
// BUFF1 162
// AND2 30
// AND3 12
// NAND4 2
// NAND3 1
// NAND8 3
// AND4 2
// NAND5 24
// AND5 16
// AND8 3
// NOR2 1

module c1908 (PNN1,PNN4,PNN7,PNN10,PNN13,PNN16,PNN19,PNN22,PNN25,PNN28,
              PNN31,PNN34,PNN37,PNN40,PNN43,PNN46,PNN49,PNN53,PNN56,PNN60,
              PNN63,PNN66,PNN69,PNN72,PNN76,PNN79,PNN82,PNN85,PNN88,PNN91,
              PNN94,PNN99,PNN104,PNN2753,PNN2754,PNN2755,PNN2756,PNN2762,PNN2767,PNN2768,
              PNN2779,PNN2780,PNN2781,PNN2782,PNN2783,PNN2784,PNN2785,PNN2786,PNN2787,PNN2811,
              PNN2886,PNN2887,PNN2888,PNN2889,PNN2890,PNN2891,PNN2892,PNN2899);

input PNN1,PNN4,PNN7,PNN10,PNN13,PNN16,PNN19,PNN22,PNN25,PNN28,
      PNN31,PNN34,PNN37,PNN40,PNN43,PNN46,PNN49,PNN53,PNN56,PNN60,
      PNN63,PNN66,PNN69,PNN72,PNN76,PNN79,PNN82,PNN85,PNN88,PNN91,
      PNN94,PNN99,PNN104;

output PNN2753,PNN2754,PNN2755,PNN2756,PNN2762,PNN2767,PNN2768,PNN2779,PNN2780,PNN2781,
       PNN2782,PNN2783,PNN2784,PNN2785,PNN2786,PNN2787,PNN2811,PNN2886,PNN2887,PNN2888,
       PNN2889,PNN2890,PNN2891,PNN2892,PNN2899;

wire PNN190,PNN194,PNN197,PNN201,PNN206,PNN209,PNN212,PNN216,PNN220,PNN225,
     PNN229,PNN232,PNN235,PNN239,PNN243,PNN247,PNN251,PNN252,PNN253,PNN256,
     PNN257,PNN260,PNN263,PNN266,PNN269,PNN272,PNN275,PNN276,PNN277,PNN280,
     PNN283,PNN290,PNN297,PNN300,PNN303,PNN306,PNN313,PNN316,PNN319,PNN326,
     PNN331,PNN338,PNN343,PNN346,PNN349,PNN352,PNN355,PNN358,PNN361,PNN364,
     PNN367,PNN370,PNN373,PNN376,PNN379,PNN382,PNN385,PNN388,PNN534,PNN535,
     PNN536,PNN537,PNN538,PNN539,PNN540,PNN541,PNN542,PNN543,PNN544,PNN545,
     PNN546,PNN547,PNN548,PNN549,PNN550,PNN551,PNN552,PNN553,PNN554,PNN555,
     PNN556,PNN559,PNN562,PNN565,PNN568,PNN571,PNN574,PNN577,PNN580,PNN583,
     PNN586,PNN589,PNN592,PNN595,PNN598,PNN601,PNN602,PNN603,PNN608,PNN612,
     PNN616,PNN619,PNN622,PNN625,PNN628,PNN631,PNN634,PNN637,PNN640,PNN643,
     PNN646,PNN649,PNN652,PNN655,PNN658,PNN661,PNN664,PNN667,PNN670,PNN673,
     PNN676,PNN679,PNN682,PNN685,PNN688,PNN691,PNN694,PNN697,PNN700,PNN703,
     PNN706,PNN709,PNN712,PNN715,PNN718,PNN721,PNN724,PNN727,PNN730,PNN733,
     PNN736,PNN739,PNN742,PNN745,PNN748,PNN751,PNN886,PNN887,PNN888,PNN889,
     PNN890,PNN891,PNN892,PNN893,PNN894,PNN895,PNN896,PNN897,PNN898,PNN899,
     PNN903,PNN907,PNN910,PNN913,PNN914,PNN915,PNN916,PNN917,PNN918,PNN919,
     PNN920,PNN921,PNN922,PNN923,PNN926,PNN935,PNN938,PNN939,PNN942,PNN943,
     PNN946,PNN947,PNN950,PNN951,PNN954,PNN955,PNN958,PNN959,PNN962,PNN965,
     PNN968,PNN969,PNN972,PNN973,PNN976,PNN977,PNN980,PNN981,PNN984,PNN985,
     PNN988,PNN989,PNN990,PNN991,PNN992,PNN993,PNN994,PNN997,PNN998,PNN1001,
     PNN1002,PNN1003,PNN1004,PNN1005,PNN1006,PNN1007,PNN1008,PNN1009,PNN1010,PNN1013,
     PNN1016,PNN1019,PNN1022,PNN1025,PNN1028,PNN1031,PNN1034,PNN1037,PNN1040,PNN1043,
     PNN1046,PNN1049,PNN1054,PNN1055,PNN1063,PNN1064,PNN1067,PNN1068,PNN1119,PNN1120,
     PNN1121,PNN1122,PNN1128,PNN1129,PNN1130,PNN1131,PNN1132,PNN1133,PNN1148,PNN1149,
     PNN1150,PNN1151,PNN1152,PNN1153,PNN1154,PNN1155,PNN1156,PNN1157,PNN1158,PNN1159,
     PNN1160,PNN1161,PNN1162,PNN1163,PNN1164,PNN1167,PNN1168,PNN1171,PNN1188,PNN1205,
     PNN1206,PNN1207,PNN1208,PNN1209,PNN1210,PNN1211,PNN1212,PNN1213,PNN1214,PNN1215,
     PNN1216,PNN1217,PNN1218,PNN1219,PNN1220,PNN1221,PNN1222,PNN1223,PNN1224,PNN1225,
     PNN1226,PNN1227,PNN1228,PNN1229,PNN1230,PNN1231,PNN1232,PNN1235,PNN1238,PNN1239,
     PNN1240,PNN1241,PNN1242,PNN1243,PNN1246,PNN1249,PNN1252,PNN1255,PNN1258,PNN1261,
     PNN1264,PNN1267,PNN1309,PNN1310,PNN1311,PNN1312,PNN1313,PNN1314,PNN1315,PNN1316,
     PNN1317,PNN1318,PNN1319,PNN1322,PNN1327,PNN1328,PNN1334,PNN1344,PNN1345,PNN1346,
     PNN1348,PNN1349,PNN1350,PNN1351,PNN1352,PNN1355,PNN1358,PNN1361,PNN1364,PNN1367,
     PNN1370,PNN1373,PNN1376,PNN1379,PNN1383,PNN1386,PNN1387,PNN1388,PNN1389,PNN1390,
     PNN1393,PNN1396,PNN1397,PNN1398,PNN1399,PNN1409,PNN1412,PNN1413,PNN1416,PNN1419,
     PNN1433,PNN1434,PNN1438,PNN1439,PNN1440,PNN1443,PNN1444,PNN1445,PNN1446,PNN1447,
     PNN1448,PNN1451,PNN1452,PNN1453,PNN1454,PNN1455,PNN1456,PNN1457,PNN1458,PNN1459,
     PNN1460,PNN1461,PNN1462,PNN1463,PNN1464,PNN1468,PNN1469,PNN1470,PNN1471,PNN1472,
     PNN1475,PNN1476,PNN1478,PNN1481,PNN1484,PNN1487,PNN1488,PNN1489,PNN1490,PNN1491,
     PNN1492,PNN1493,PNN1494,PNN1495,PNN1496,PNN1498,PNN1499,PNN1500,PNN1501,PNN1504,
     PNN1510,PNN1513,PNN1514,PNN1517,PNN1520,PNN1521,PNN1522,PNN1526,PNN1527,PNN1528,
     PNN1529,PNN1530,PNN1531,PNN1532,PNN1534,PNN1537,PNN1540,PNN1546,PNN1554,PNN1557,
     PNN1561,PNN1567,PNN1568,PNN1569,PNN1571,PNN1576,PNN1588,PNN1591,PNN1593,PNN1594,
     PNN1595,PNN1596,PNN1600,PNN1603,PNN1606,PNN1609,PNN1612,PNN1615,PNN1620,PNN1623,
     PNN1635,PNN1636,PNN1638,PNN1639,PNN1640,PNN1643,PNN1647,PNN1651,PNN1658,PNN1661,
     PNN1664,PNN1671,PNN1672,PNN1675,PNN1677,PNN1678,PNN1679,PNN1680,PNN1681,PNN1682,
     PNN1683,PNN1685,PNN1688,PNN1697,PNN1701,PNN1706,PNN1707,PNN1708,PNN1709,PNN1710,
     PNN1711,PNN1712,PNN1713,PNN1714,PNN1717,PNN1720,PNN1721,PNN1723,PNN1727,PNN1728,
     PNN1730,PNN1731,PNN1734,PNN1740,PNN1741,PNN1742,PNN1746,PNN1747,PNN1748,PNN1751,
     PNN1759,PNN1761,PNN1762,PNN1763,PNN1764,PNN1768,PNN1769,PNN1772,PNN1773,PNN1774,
     PNN1777,PNN1783,PNN1784,PNN1785,PNN1786,PNN1787,PNN1788,PNN1791,PNN1792,PNN1795,
     PNN1796,PNN1798,PNN1801,PNN1802,PNN1807,PNN1808,PNN1809,PNN1810,PNN1812,PNN1815,
     PNN1818,PNN1821,PNN1822,PNN1823,PNN1824,PNN1825,PNN1826,PNN1827,PNN1830,PNN1837,
     PNN1838,PNN1841,PNN1848,PNN1849,PNN1850,PNN1852,PNN1855,PNN1856,PNN1857,PNN1858,
     PNN1864,PNN1865,PNN1866,PNN1869,PNN1872,PNN1875,PNN1878,PNN1879,PNN1882,PNN1883,
     PNN1884,PNN1885,PNN1889,PNN1895,PNN1896,PNN1897,PNN1898,PNN1902,PNN1910,PNN1911,
     PNN1912,PNN1913,PNN1915,PNN1919,PNN1920,PNN1921,PNN1922,PNN1923,PNN1924,PNN1927,
     PNN1930,PNN1933,PNN1936,PNN1937,PNN1938,PNN1941,PNN1942,PNN1944,PNN1947,PNN1950,
     PNN1953,PNN1958,PNN1961,PNN1965,PNN1968,PNN1975,PNN1976,PNN1977,PNN1978,PNN1979,
     PNN1980,PNN1985,PNN1987,PNN1999,PNN2000,PNN2002,PNN2003,PNN2004,PNN2005,PNN2006,
     PNN2007,PNN2008,PNN2009,PNN2012,PNN2013,PNN2014,PNN2015,PNN2016,PNN2018,PNN2019,
     PNN2020,PNN2021,PNN2022,PNN2023,PNN2024,PNN2025,PNN2026,PNN2027,PNN2030,PNN2033,
     PNN2036,PNN2037,PNN2038,PNN2039,PNN2040,PNN2041,PNN2042,PNN2047,PNN2052,PNN2055,
     PNN2060,PNN2061,PNN2062,PNN2067,PNN2068,PNN2071,PNN2076,PNN2077,PNN2078,PNN2081,
     PNN2086,PNN2089,PNN2104,PNN2119,PNN2129,PNN2143,PNN2148,PNN2151,PNN2196,PNN2199,
     PNN2202,PNN2205,PNN2214,PNN2215,PNN2216,PNN2217,PNN2222,PNN2223,PNN2224,PNN2225,
     PNN2226,PNN2227,PNN2228,PNN2229,PNN2230,PNN2231,PNN2232,PNN2233,PNN2234,PNN2235,
     PNN2236,PNN2237,PNN2240,PNN2241,PNN2244,PNN2245,PNN2250,PNN2253,PNN2256,PNN2257,
     PNN2260,PNN2263,PNN2266,PNN2269,PNN2272,PNN2279,PNN2286,PNN2297,PNN2315,PNN2326,
     PNN2340,PNN2353,PNN2361,PNN2375,PNN2384,PNN2385,PNN2386,PNN2426,PNN2427,PNN2537,
     PNN2540,PNN2543,PNN2546,PNN2549,PNN2552,PNN2555,PNN2558,PNN2561,PNN2564,PNN2567,
     PNN2570,PNN2573,PNN2576,PNN2594,PNN2597,PNN2600,PNN2603,PNN2606,PNN2611,PNN2614,
     PNN2617,PNN2620,PNN2627,PNN2628,PNN2629,PNN2630,PNN2631,PNN2632,PNN2633,PNN2634,
     PNN2639,PNN2642,PNN2645,PNN2648,PNN2651,PNN2655,PNN2658,PNN2661,PNN2664,PNN2669,
     PNN2670,PNN2671,PNN2672,PNN2673,PNN2674,PNN2675,PNN2676,PNN2682,PNN2683,PNN2688,
     PNN2689,PNN2690,PNN2691,PNN2710,PNN2720,PNN2721,PNN2722,PNN2723,PNN2724,PNN2725,
     PNN2726,PNN2727,PNN2728,PNN2729,PNN2730,PNN2731,PNN2732,PNN2733,PNN2734,PNN2735,
     PNN2736,PNN2737,PNN2738,PNN2739,PNN2740,PNN2741,PNN2742,PNN2743,PNN2744,PNN2745,
     PNN2746,PNN2747,PNN2750,PNN2757,PNN2758,PNN2759,PNN2760,PNN2761,PNN2763,PNN2764,
     PNN2765,PNN2766,PNN2773,PNN2776,PNN2788,PNN2789,PNN2800,PNN2807,PNN2808,PNN2809,
     PNN2810,PNN2812,PNN2815,PNN2818,PNN2821,PNN2824,PNN2827,PNN2828,PNN2829,PNN2843,
     PNN2846,PNN2850,PNN2851,PNN2852,PNN2853,PNN2854,PNN2857,PNN2858,PNN2859,PNN2860,
     PNN2861,PNN2862,PNN2863,PNN2866,PNN2867,PNN2868,PNN2869,PNN2870,PNN2871,PNN2872,
     PNN2873,PNN2874,PNN2875,PNN2876,PNN2877,PNN2878,PNN2879,PNN2880,PNN2881,PNN2882,
     PNN2883,PNN2895,PNN2896,PNN2897,PNN2898;

not NOT1_1 (PNN190, PNN1);
not NOT1_2 (PNN194, PNN4);
not NOT1_3 (PNN197, PNN7);
not NOT1_4 (PNN201, PNN10);
not NOT1_5 (PNN206, PNN13);
not NOT1_6 (PNN209, PNN16);
not NOT1_7 (PNN212, PNN19);
not NOT1_8 (PNN216, PNN22);
not NOT1_9 (PNN220, PNN25);
not NOT1_10 (PNN225, PNN28);
not NOT1_11 (PNN229, PNN31);
not NOT1_12 (PNN232, PNN34);
not NOT1_13 (PNN235, PNN37);
not NOT1_14 (PNN239, PNN40);
not NOT1_15 (PNN243, PNN43);
not NOT1_16 (PNN247, PNN46);
nand NAND2_17 (PNN251, PNN63, PNN88);
nand NAND2_18 (PNN252, PNN66, PNN91);
not NOT1_19 (PNN253, PNN72);
not NOT1_20 (PNN256, PNN72);
buf BUFF1_21 (PNN257, PNN69);
buf BUFF1_22 (PNN260, PNN69);
not NOT1_23 (PNN263, PNN76);
not NOT1_24 (PNN266, PNN79);
not NOT1_25 (PNN269, PNN82);
not NOT1_26 (PNN272, PNN85);
not NOT1_27 (PNN275, PNN104);
not NOT1_28 (PNN276, PNN104);
not NOT1_29 (PNN277, PNN88);
not NOT1_30 (PNN280, PNN91);
buf BUFF1_31 (PNN283, PNN94);
not NOT1_32 (PNN290, PNN94);
buf BUFF1_33 (PNN297, PNN94);
not NOT1_34 (PNN300, PNN94);
buf BUFF1_35 (PNN303, PNN99);
not NOT1_36 (PNN306, PNN99);
not NOT1_37 (PNN313, PNN99);
buf BUFF1_38 (PNN316, PNN104);
not NOT1_39 (PNN319, PNN104);
buf BUFF1_40 (PNN326, PNN104);
buf BUFF1_41 (PNN331, PNN104);
not NOT1_42 (PNN338, PNN104);
buf BUFF1_43 (PNN343, PNN1);
buf BUFF1_44 (PNN346, PNN4);
buf BUFF1_45 (PNN349, PNN7);
buf BUFF1_46 (PNN352, PNN10);
buf BUFF1_47 (PNN355, PNN13);
buf BUFF1_48 (PNN358, PNN16);
buf BUFF1_49 (PNN361, PNN19);
buf BUFF1_50 (PNN364, PNN22);
buf BUFF1_51 (PNN367, PNN25);
buf BUFF1_52 (PNN370, PNN28);
buf BUFF1_53 (PNN373, PNN31);
buf BUFF1_54 (PNN376, PNN34);
buf BUFF1_55 (PNN379, PNN37);
buf BUFF1_56 (PNN382, PNN40);
buf BUFF1_57 (PNN385, PNN43);
buf BUFF1_58 (PNN388, PNN46);
not NOT1_59 (PNN534, PNN343);
not NOT1_60 (PNN535, PNN346);
not NOT1_61 (PNN536, PNN349);
not NOT1_62 (PNN537, PNN352);
not NOT1_63 (PNN538, PNN355);
not NOT1_64 (PNN539, PNN358);
not NOT1_65 (PNN540, PNN361);
not NOT1_66 (PNN541, PNN364);
not NOT1_67 (PNN542, PNN367);
not NOT1_68 (PNN543, PNN370);
not NOT1_69 (PNN544, PNN373);
not NOT1_70 (PNN545, PNN376);
not NOT1_71 (PNN546, PNN379);
not NOT1_72 (PNN547, PNN382);
not NOT1_73 (PNN548, PNN385);
not NOT1_74 (PNN549, PNN388);
nand NAND2_75 (PNN550, PNN306, PNN331);
nand NAND2_76 (PNN551, PNN306, PNN331);
nand NAND2_77 (PNN552, PNN306, PNN331);
nand NAND2_78 (PNN553, PNN306, PNN331);
nand NAND2_79 (PNN554, PNN306, PNN331);
nand NAND2_80 (PNN555, PNN306, PNN331);
buf BUFF1_81 (PNN556, PNN190);
buf BUFF1_82 (PNN559, PNN194);
buf BUFF1_83 (PNN562, PNN206);
buf BUFF1_84 (PNN565, PNN209);
buf BUFF1_85 (PNN568, PNN225);
buf BUFF1_86 (PNN571, PNN243);
and AND2_87 (PNN574, PNN63, PNN319);
buf BUFF1_88 (PNN577, PNN220);
buf BUFF1_89 (PNN580, PNN229);
buf BUFF1_90 (PNN583, PNN232);
and AND2_91 (PNN586, PNN66, PNN319);
buf BUFF1_92 (PNN589, PNN239);
and AND3_93 (PNN592, PNN49, PNN253, PNN319);
buf BUFF1_94 (PNN595, PNN247);
buf BUFF1_95 (PNN598, PNN239);
nand NAND2_96 (PNN601, PNN326, PNN277);
nand NAND2_97 (PNN602, PNN326, PNN280);
nand NAND2_98 (PNN603, PNN260, PNN72);
nand NAND2_99 (PNN608, PNN260, PNN300);
nand NAND2_100 (PNN612, PNN256, PNN300);
buf BUFF1_101 (PNN616, PNN201);
buf BUFF1_102 (PNN619, PNN216);
buf BUFF1_103 (PNN622, PNN220);
buf BUFF1_104 (PNN625, PNN239);
buf BUFF1_105 (PNN628, PNN190);
buf BUFF1_106 (PNN631, PNN190);
buf BUFF1_107 (PNN634, PNN194);
buf BUFF1_108 (PNN637, PNN229);
buf BUFF1_109 (PNN640, PNN197);
and AND3_110 (PNN643, PNN56, PNN257, PNN319);
buf BUFF1_111 (PNN646, PNN232);
buf BUFF1_112 (PNN649, PNN201);
buf BUFF1_113 (PNN652, PNN235);
and AND3_114 (PNN655, PNN60, PNN257, PNN319);
buf BUFF1_115 (PNN658, PNN263);
buf BUFF1_116 (PNN661, PNN263);
buf BUFF1_117 (PNN664, PNN266);
buf BUFF1_118 (PNN667, PNN266);
buf BUFF1_119 (PNN670, PNN269);
buf BUFF1_120 (PNN673, PNN269);
buf BUFF1_121 (PNN676, PNN272);
buf BUFF1_122 (PNN679, PNN272);
and AND2_123 (PNN682, PNN251, PNN316);
and AND2_124 (PNN685, PNN252, PNN316);
buf BUFF1_125 (PNN688, PNN197);
buf BUFF1_126 (PNN691, PNN197);
buf BUFF1_127 (PNN694, PNN212);
buf BUFF1_128 (PNN697, PNN212);
buf BUFF1_129 (PNN700, PNN247);
buf BUFF1_130 (PNN703, PNN247);
buf BUFF1_131 (PNN706, PNN235);
buf BUFF1_132 (PNN709, PNN235);
buf BUFF1_133 (PNN712, PNN201);
buf BUFF1_134 (PNN715, PNN201);
buf BUFF1_135 (PNN718, PNN206);
buf BUFF1_136 (PNN721, PNN216);
and AND3_137 (PNN724, PNN53, PNN253, PNN319);
buf BUFF1_138 (PNN727, PNN243);
buf BUFF1_139 (PNN730, PNN220);
buf BUFF1_140 (PNN733, PNN220);
buf BUFF1_141 (PNN736, PNN209);
buf BUFF1_142 (PNN739, PNN216);
buf BUFF1_143 (PNN742, PNN225);
buf BUFF1_144 (PNN745, PNN243);
buf BUFF1_145 (PNN748, PNN212);
buf BUFF1_146 (PNN751, PNN225);
not NOT1_147 (PNN886, PNN682);
not NOT1_148 (PNN887, PNN685);
not NOT1_149 (PNN888, PNN616);
not NOT1_150 (PNN889, PNN619);
not NOT1_151 (PNN890, PNN622);
not NOT1_152 (PNN891, PNN625);
not NOT1_153 (PNN892, PNN631);
not NOT1_154 (PNN893, PNN643);
not NOT1_155 (PNN894, PNN649);
not NOT1_156 (PNN895, PNN652);
not NOT1_157 (PNN896, PNN655);
and AND2_158 (PNN897, PNN49, PNN612);
and AND2_159 (PNN898, PNN56, PNN608);
nand NAND2_160 (PNN899, PNN53, PNN612);
nand NAND2_161 (PNN903, PNN60, PNN608);
nand NAND2_162 (PNN907, PNN49, PNN612);
nand NAND2_163 (PNN910, PNN56, PNN608);
not NOT1_164 (PNN913, PNN661);
not NOT1_165 (PNN914, PNN658);
not NOT1_166 (PNN915, PNN667);
not NOT1_167 (PNN916, PNN664);
not NOT1_168 (PNN917, PNN673);
not NOT1_169 (PNN918, PNN670);
not NOT1_170 (PNN919, PNN679);
not NOT1_171 (PNN920, PNN676);
nand NAND4_172 (PNN921, PNN277, PNN297, PNN326, PNN603);
nand NAND4_173 (PNN922, PNN280, PNN297, PNN326, PNN603);
nand NAND3_174 (PNN923, PNN303, PNN338, PNN603);
and AND3_175 (PNN926, PNN303, PNN338, PNN603);
buf BUFF1_176 (PNN935, PNN556);
not NOT1_177 (PNN938, PNN688);
buf BUFF1_178 (PNN939, PNN556);
not NOT1_179 (PNN942, PNN691);
buf BUFF1_180 (PNN943, PNN562);
not NOT1_181 (PNN946, PNN694);
buf BUFF1_182 (PNN947, PNN562);
not NOT1_183 (PNN950, PNN697);
buf BUFF1_184 (PNN951, PNN568);
not NOT1_185 (PNN954, PNN700);
buf BUFF1_186 (PNN955, PNN568);
not NOT1_187 (PNN958, PNN703);
buf BUFF1_188 (PNN959, PNN574);
buf BUFF1_189 (PNN962, PNN574);
buf BUFF1_190 (PNN965, PNN580);
not NOT1_191 (PNN968, PNN706);
buf BUFF1_192 (PNN969, PNN580);
not NOT1_193 (PNN972, PNN709);
buf BUFF1_194 (PNN973, PNN586);
not NOT1_195 (PNN976, PNN712);
buf BUFF1_196 (PNN977, PNN586);
not NOT1_197 (PNN980, PNN715);
buf BUFF1_198 (PNN981, PNN592);
not NOT1_199 (PNN984, PNN628);
buf BUFF1_200 (PNN985, PNN592);
not NOT1_201 (PNN988, PNN718);
not NOT1_202 (PNN989, PNN721);
not NOT1_203 (PNN990, PNN634);
not NOT1_204 (PNN991, PNN724);
not NOT1_205 (PNN992, PNN727);
not NOT1_206 (PNN993, PNN637);
buf BUFF1_207 (PNN994, PNN595);
not NOT1_208 (PNN997, PNN730);
buf BUFF1_209 (PNN998, PNN595);
not NOT1_210 (PNN1001, PNN733);
not NOT1_211 (PNN1002, PNN736);
not NOT1_212 (PNN1003, PNN739);
not NOT1_213 (PNN1004, PNN640);
not NOT1_214 (PNN1005, PNN742);
not NOT1_215 (PNN1006, PNN745);
not NOT1_216 (PNN1007, PNN646);
not NOT1_217 (PNN1008, PNN748);
not NOT1_218 (PNN1009, PNN751);
buf BUFF1_219 (PNN1010, PNN559);
buf BUFF1_220 (PNN1013, PNN559);
buf BUFF1_221 (PNN1016, PNN565);
buf BUFF1_222 (PNN1019, PNN565);
buf BUFF1_223 (PNN1022, PNN571);
buf BUFF1_224 (PNN1025, PNN571);
buf BUFF1_225 (PNN1028, PNN577);
buf BUFF1_226 (PNN1031, PNN577);
buf BUFF1_227 (PNN1034, PNN583);
buf BUFF1_228 (PNN1037, PNN583);
buf BUFF1_229 (PNN1040, PNN589);
buf BUFF1_230 (PNN1043, PNN589);
buf BUFF1_231 (PNN1046, PNN598);
buf BUFF1_232 (PNN1049, PNN598);
nand NAND2_233 (PNN1054, PNN619, PNN888);
nand NAND2_234 (PNN1055, PNN616, PNN889);
nand NAND2_235 (PNN1063, PNN625, PNN890);
nand NAND2_236 (PNN1064, PNN622, PNN891);
nand NAND2_237 (PNN1067, PNN655, PNN895);
nand NAND2_238 (PNN1068, PNN652, PNN896);
nand NAND2_239 (PNN1119, PNN721, PNN988);
nand NAND2_240 (PNN1120, PNN718, PNN989);
nand NAND2_241 (PNN1121, PNN727, PNN991);
nand NAND2_242 (PNN1122, PNN724, PNN992);
nand NAND2_243 (PNN1128, PNN739, PNN1002);
nand NAND2_244 (PNN1129, PNN736, PNN1003);
nand NAND2_245 (PNN1130, PNN745, PNN1005);
nand NAND2_246 (PNN1131, PNN742, PNN1006);
nand NAND2_247 (PNN1132, PNN751, PNN1008);
nand NAND2_248 (PNN1133, PNN748, PNN1009);
not NOT1_249 (PNN1148, PNN939);
not NOT1_250 (PNN1149, PNN935);
nand NAND2_251 (PNN1150, PNN1054, PNN1055);
not NOT1_252 (PNN1151, PNN943);
not NOT1_253 (PNN1152, PNN947);
not NOT1_254 (PNN1153, PNN955);
not NOT1_255 (PNN1154, PNN951);
not NOT1_256 (PNN1155, PNN962);
not NOT1_257 (PNN1156, PNN969);
not NOT1_258 (PNN1157, PNN977);
nand NAND2_259 (PNN1158, PNN1063, PNN1064);
not NOT1_260 (PNN1159, PNN985);
nand NAND2_261 (PNN1160, PNN985, PNN892);
not NOT1_262 (PNN1161, PNN998);
nand NAND2_263 (PNN1162, PNN1067, PNN1068);
not NOT1_264 (PNN1163, PNN899);
buf BUFF1_265 (PNN1164, PNN899);
not NOT1_266 (PNN1167, PNN903);
buf BUFF1_267 (PNN1168, PNN903);
nand NAND2_268 (PNN1171, PNN921, PNN923);
nand NAND2_269 (PNN1188, PNN922, PNN923);
not NOT1_270 (PNN1205, PNN1010);
nand NAND2_271 (PNN1206, PNN1010, PNN938);
not NOT1_272 (PNN1207, PNN1013);
nand NAND2_273 (PNN1208, PNN1013, PNN942);
not NOT1_274 (PNN1209, PNN1016);
nand NAND2_275 (PNN1210, PNN1016, PNN946);
not NOT1_276 (PNN1211, PNN1019);
nand NAND2_277 (PNN1212, PNN1019, PNN950);
not NOT1_278 (PNN1213, PNN1022);
nand NAND2_279 (PNN1214, PNN1022, PNN954);
not NOT1_280 (PNN1215, PNN1025);
nand NAND2_281 (PNN1216, PNN1025, PNN958);
not NOT1_282 (PNN1217, PNN1028);
not NOT1_283 (PNN1218, PNN959);
not NOT1_284 (PNN1219, PNN1031);
not NOT1_285 (PNN1220, PNN1034);
nand NAND2_286 (PNN1221, PNN1034, PNN968);
not NOT1_287 (PNN1222, PNN965);
not NOT1_288 (PNN1223, PNN1037);
nand NAND2_289 (PNN1224, PNN1037, PNN972);
not NOT1_290 (PNN1225, PNN1040);
nand NAND2_291 (PNN1226, PNN1040, PNN976);
not NOT1_292 (PNN1227, PNN973);
not NOT1_293 (PNN1228, PNN1043);
nand NAND2_294 (PNN1229, PNN1043, PNN980);
not NOT1_295 (PNN1230, PNN981);
nand NAND2_296 (PNN1231, PNN981, PNN984);
nand NAND2_297 (PNN1232, PNN1119, PNN1120);
nand NAND2_298 (PNN1235, PNN1121, PNN1122);
not NOT1_299 (PNN1238, PNN1046);
nand NAND2_300 (PNN1239, PNN1046, PNN997);
not NOT1_301 (PNN1240, PNN994);
not NOT1_302 (PNN1241, PNN1049);
nand NAND2_303 (PNN1242, PNN1049, PNN1001);
nand NAND2_304 (PNN1243, PNN1128, PNN1129);
nand NAND2_305 (PNN1246, PNN1130, PNN1131);
nand NAND2_306 (PNN1249, PNN1132, PNN1133);
buf BUFF1_307 (PNN1252, PNN907);
buf BUFF1_308 (PNN1255, PNN907);
buf BUFF1_309 (PNN1258, PNN910);
buf BUFF1_310 (PNN1261, PNN910);
not NOT1_311 (PNN1264, PNN1150);
nand NAND2_312 (PNN1267, PNN631, PNN1159);
nand NAND2_313 (PNN1309, PNN688, PNN1205);
nand NAND2_314 (PNN1310, PNN691, PNN1207);
nand NAND2_315 (PNN1311, PNN694, PNN1209);
nand NAND2_316 (PNN1312, PNN697, PNN1211);
nand NAND2_317 (PNN1313, PNN700, PNN1213);
nand NAND2_318 (PNN1314, PNN703, PNN1215);
nand NAND2_319 (PNN1315, PNN706, PNN1220);
nand NAND2_320 (PNN1316, PNN709, PNN1223);
nand NAND2_321 (PNN1317, PNN712, PNN1225);
nand NAND2_322 (PNN1318, PNN715, PNN1228);
not NOT1_323 (PNN1319, PNN1158);
nand NAND2_324 (PNN1322, PNN628, PNN1230);
nand NAND2_325 (PNN1327, PNN730, PNN1238);
nand NAND2_326 (PNN1328, PNN733, PNN1241);
not NOT1_327 (PNN1334, PNN1162);
nand NAND2_328 (PNN1344, PNN1267, PNN1160);
nand NAND2_329 (PNN1345, PNN1249, PNN894);
not NOT1_330 (PNN1346, PNN1249);
not NOT1_331 (PNN1348, PNN1255);
not NOT1_332 (PNN1349, PNN1252);
not NOT1_333 (PNN1350, PNN1261);
not NOT1_334 (PNN1351, PNN1258);
nand NAND2_335 (PNN1352, PNN1309, PNN1206);
nand NAND2_336 (PNN1355, PNN1310, PNN1208);
nand NAND2_337 (PNN1358, PNN1311, PNN1210);
nand NAND2_338 (PNN1361, PNN1312, PNN1212);
nand NAND2_339 (PNN1364, PNN1313, PNN1214);
nand NAND2_340 (PNN1367, PNN1314, PNN1216);
nand NAND2_341 (PNN1370, PNN1315, PNN1221);
nand NAND2_342 (PNN1373, PNN1316, PNN1224);
nand NAND2_343 (PNN1376, PNN1317, PNN1226);
nand NAND2_344 (PNN1379, PNN1318, PNN1229);
nand NAND2_345 (PNN1383, PNN1322, PNN1231);
not NOT1_346 (PNN1386, PNN1232);
nand NAND2_347 (PNN1387, PNN1232, PNN990);
not NOT1_348 (PNN1388, PNN1235);
nand NAND2_349 (PNN1389, PNN1235, PNN993);
nand NAND2_350 (PNN1390, PNN1327, PNN1239);
nand NAND2_351 (PNN1393, PNN1328, PNN1242);
not NOT1_352 (PNN1396, PNN1243);
nand NAND2_353 (PNN1397, PNN1243, PNN1004);
not NOT1_354 (PNN1398, PNN1246);
nand NAND2_355 (PNN1399, PNN1246, PNN1007);
not NOT1_356 (PNN1409, PNN1319);
nand NAND2_357 (PNN1412, PNN649, PNN1346);
not NOT1_358 (PNN1413, PNN1334);
buf BUFF1_359 (PNN1416, PNN1264);
buf BUFF1_360 (PNN1419, PNN1264);
nand NAND2_361 (PNN1433, PNN634, PNN1386);
nand NAND2_362 (PNN1434, PNN637, PNN1388);
nand NAND2_363 (PNN1438, PNN640, PNN1396);
nand NAND2_364 (PNN1439, PNN646, PNN1398);
not NOT1_365 (PNN1440, PNN1344);
nand NAND2_366 (PNN1443, PNN1355, PNN1148);
not NOT1_367 (PNN1444, PNN1355);
nand NAND2_368 (PNN1445, PNN1352, PNN1149);
not NOT1_369 (PNN1446, PNN1352);
nand NAND2_370 (PNN1447, PNN1358, PNN1151);
not NOT1_371 (PNN1448, PNN1358);
nand NAND2_372 (PNN1451, PNN1361, PNN1152);
not NOT1_373 (PNN1452, PNN1361);
nand NAND2_374 (PNN1453, PNN1367, PNN1153);
not NOT1_375 (PNN1454, PNN1367);
nand NAND2_376 (PNN1455, PNN1364, PNN1154);
not NOT1_377 (PNN1456, PNN1364);
nand NAND2_378 (PNN1457, PNN1373, PNN1156);
not NOT1_379 (PNN1458, PNN1373);
nand NAND2_380 (PNN1459, PNN1379, PNN1157);
not NOT1_381 (PNN1460, PNN1379);
not NOT1_382 (PNN1461, PNN1383);
nand NAND2_383 (PNN1462, PNN1393, PNN1161);
not NOT1_384 (PNN1463, PNN1393);
nand NAND2_385 (PNN1464, PNN1345, PNN1412);
not NOT1_386 (PNN1468, PNN1370);
nand NAND2_387 (PNN1469, PNN1370, PNN1222);
not NOT1_388 (PNN1470, PNN1376);
nand NAND2_389 (PNN1471, PNN1376, PNN1227);
nand NAND2_390 (PNN1472, PNN1387, PNN1433);
not NOT1_391 (PNN1475, PNN1390);
nand NAND2_392 (PNN1476, PNN1390, PNN1240);
nand NAND2_393 (PNN1478, PNN1389, PNN1434);
nand NAND2_394 (PNN1481, PNN1399, PNN1439);
nand NAND2_395 (PNN1484, PNN1397, PNN1438);
nand NAND2_396 (PNN1487, PNN939, PNN1444);
nand NAND2_397 (PNN1488, PNN935, PNN1446);
nand NAND2_398 (PNN1489, PNN943, PNN1448);
not NOT1_399 (PNN1490, PNN1419);
not NOT1_400 (PNN1491, PNN1416);
nand NAND2_401 (PNN1492, PNN947, PNN1452);
nand NAND2_402 (PNN1493, PNN955, PNN1454);
nand NAND2_403 (PNN1494, PNN951, PNN1456);
nand NAND2_404 (PNN1495, PNN969, PNN1458);
nand NAND2_405 (PNN1496, PNN977, PNN1460);
nand NAND2_406 (PNN1498, PNN998, PNN1463);
not NOT1_407 (PNN1499, PNN1440);
nand NAND2_408 (PNN1500, PNN965, PNN1468);
nand NAND2_409 (PNN1501, PNN973, PNN1470);
nand NAND2_410 (PNN1504, PNN994, PNN1475);
not NOT1_411 (PNN1510, PNN1464);
nand NAND2_412 (PNN1513, PNN1443, PNN1487);
nand NAND2_413 (PNN1514, PNN1445, PNN1488);
nand NAND2_414 (PNN1517, PNN1447, PNN1489);
nand NAND2_415 (PNN1520, PNN1451, PNN1492);
nand NAND2_416 (PNN1521, PNN1453, PNN1493);
nand NAND2_417 (PNN1522, PNN1455, PNN1494);
nand NAND2_418 (PNN1526, PNN1457, PNN1495);
nand NAND2_419 (PNN1527, PNN1459, PNN1496);
not NOT1_420 (PNN1528, PNN1472);
nand NAND2_421 (PNN1529, PNN1462, PNN1498);
not NOT1_422 (PNN1530, PNN1478);
not NOT1_423 (PNN1531, PNN1481);
not NOT1_424 (PNN1532, PNN1484);
nand NAND2_425 (PNN1534, PNN1471, PNN1501);
nand NAND2_426 (PNN1537, PNN1469, PNN1500);
nand NAND2_427 (PNN1540, PNN1476, PNN1504);
not NOT1_428 (PNN1546, PNN1513);
not NOT1_429 (PNN1554, PNN1521);
not NOT1_430 (PNN1557, PNN1526);
not NOT1_431 (PNN1561, PNN1520);
nand NAND2_432 (PNN1567, PNN1484, PNN1531);
nand NAND2_433 (PNN1568, PNN1481, PNN1532);
not NOT1_434 (PNN1569, PNN1510);
not NOT1_435 (PNN1571, PNN1527);
not NOT1_436 (PNN1576, PNN1529);
buf BUFF1_437 (PNN1588, PNN1522);
not NOT1_438 (PNN1591, PNN1534);
not NOT1_439 (PNN1593, PNN1537);
nand NAND2_440 (PNN1594, PNN1540, PNN1530);
not NOT1_441 (PNN1595, PNN1540);
nand NAND2_442 (PNN1596, PNN1567, PNN1568);
buf BUFF1_443 (PNN1600, PNN1517);
buf BUFF1_444 (PNN1603, PNN1517);
buf BUFF1_445 (PNN1606, PNN1522);
buf BUFF1_446 (PNN1609, PNN1522);
buf BUFF1_447 (PNN1612, PNN1514);
buf BUFF1_448 (PNN1615, PNN1514);
buf BUFF1_449 (PNN1620, PNN1557);
buf BUFF1_450 (PNN1623, PNN1554);
not NOT1_451 (PNN1635, PNN1571);
nand NAND2_452 (PNN1636, PNN1478, PNN1595);
nand NAND2_453 (PNN1638, PNN1576, PNN1569);
not NOT1_454 (PNN1639, PNN1576);
buf BUFF1_455 (PNN1640, PNN1561);
buf BUFF1_456 (PNN1643, PNN1561);
buf BUFF1_457 (PNN1647, PNN1546);
buf BUFF1_458 (PNN1651, PNN1546);
buf BUFF1_459 (PNN1658, PNN1554);
buf BUFF1_460 (PNN1661, PNN1557);
buf BUFF1_461 (PNN1664, PNN1557);
nand NAND2_462 (PNN1671, PNN1596, PNN893);
not NOT1_463 (PNN1672, PNN1596);
not NOT1_464 (PNN1675, PNN1600);
not NOT1_465 (PNN1677, PNN1603);
nand NAND2_466 (PNN1678, PNN1606, PNN1217);
not NOT1_467 (PNN1679, PNN1606);
nand NAND2_468 (PNN1680, PNN1609, PNN1219);
not NOT1_469 (PNN1681, PNN1609);
not NOT1_470 (PNN1682, PNN1612);
not NOT1_471 (PNN1683, PNN1615);
nand NAND2_472 (PNN1685, PNN1594, PNN1636);
nand NAND2_473 (PNN1688, PNN1510, PNN1639);
buf BUFF1_474 (PNN1697, PNN1588);
buf BUFF1_475 (PNN1701, PNN1588);
nand NAND2_476 (PNN1706, PNN643, PNN1672);
not NOT1_477 (PNN1707, PNN1643);
nand NAND2_478 (PNN1708, PNN1647, PNN1675);
not NOT1_479 (PNN1709, PNN1647);
nand NAND2_480 (PNN1710, PNN1651, PNN1677);
not NOT1_481 (PNN1711, PNN1651);
nand NAND2_482 (PNN1712, PNN1028, PNN1679);
nand NAND2_483 (PNN1713, PNN1031, PNN1681);
buf BUFF1_484 (PNN1714, PNN1620);
buf BUFF1_485 (PNN1717, PNN1620);
nand NAND2_486 (PNN1720, PNN1658, PNN1593);
not NOT1_487 (PNN1721, PNN1658);
nand NAND2_488 (PNN1723, PNN1638, PNN1688);
not NOT1_489 (PNN1727, PNN1661);
not NOT1_490 (PNN1728, PNN1640);
not NOT1_491 (PNN1730, PNN1664);
buf BUFF1_492 (PNN1731, PNN1623);
buf BUFF1_493 (PNN1734, PNN1623);
nand NAND2_494 (PNN1740, PNN1685, PNN1528);
not NOT1_495 (PNN1741, PNN1685);
nand NAND2_496 (PNN1742, PNN1671, PNN1706);
nand NAND2_497 (PNN1746, PNN1600, PNN1709);
nand NAND2_498 (PNN1747, PNN1603, PNN1711);
nand NAND2_499 (PNN1748, PNN1678, PNN1712);
nand NAND2_500 (PNN1751, PNN1680, PNN1713);
nand NAND2_501 (PNN1759, PNN1537, PNN1721);
not NOT1_502 (PNN1761, PNN1697);
nand NAND2_503 (PNN1762, PNN1697, PNN1727);
not NOT1_504 (PNN1763, PNN1701);
nand NAND2_505 (PNN1764, PNN1701, PNN1730);
not NOT1_506 (PNN1768, PNN1717);
nand NAND2_507 (PNN1769, PNN1472, PNN1741);
nand NAND2_508 (PNN1772, PNN1723, PNN1413);
not NOT1_509 (PNN1773, PNN1723);
nand NAND2_510 (PNN1774, PNN1708, PNN1746);
nand NAND2_511 (PNN1777, PNN1710, PNN1747);
not NOT1_512 (PNN1783, PNN1731);
nand NAND2_513 (PNN1784, PNN1731, PNN1682);
not NOT1_514 (PNN1785, PNN1714);
not NOT1_515 (PNN1786, PNN1734);
nand NAND2_516 (PNN1787, PNN1734, PNN1683);
nand NAND2_517 (PNN1788, PNN1720, PNN1759);
nand NAND2_518 (PNN1791, PNN1661, PNN1761);
nand NAND2_519 (PNN1792, PNN1664, PNN1763);
nand NAND2_520 (PNN1795, PNN1751, PNN1155);
not NOT1_521 (PNN1796, PNN1751);
nand NAND2_522 (PNN1798, PNN1740, PNN1769);
nand NAND2_523 (PNN1801, PNN1334, PNN1773);
nand NAND2_524 (PNN1802, PNN1742, PNN290);
not NOT1_525 (PNN1807, PNN1748);
nand NAND2_526 (PNN1808, PNN1748, PNN1218);
nand NAND2_527 (PNN1809, PNN1612, PNN1783);
nand NAND2_528 (PNN1810, PNN1615, PNN1786);
nand NAND2_529 (PNN1812, PNN1791, PNN1762);
nand NAND2_530 (PNN1815, PNN1792, PNN1764);
buf BUFF1_531 (PNN1818, PNN1742);
nand NAND2_532 (PNN1821, PNN1777, PNN1490);
not NOT1_533 (PNN1822, PNN1777);
nand NAND2_534 (PNN1823, PNN1774, PNN1491);
not NOT1_535 (PNN1824, PNN1774);
nand NAND2_536 (PNN1825, PNN962, PNN1796);
nand NAND2_537 (PNN1826, PNN1788, PNN1409);
not NOT1_538 (PNN1827, PNN1788);
nand NAND2_539 (PNN1830, PNN1772, PNN1801);
nand NAND2_540 (PNN1837, PNN959, PNN1807);
nand NAND2_541 (PNN1838, PNN1809, PNN1784);
nand NAND2_542 (PNN1841, PNN1810, PNN1787);
nand NAND2_543 (PNN1848, PNN1419, PNN1822);
nand NAND2_544 (PNN1849, PNN1416, PNN1824);
nand NAND2_545 (PNN1850, PNN1795, PNN1825);
nand NAND2_546 (PNN1852, PNN1319, PNN1827);
nand NAND2_547 (PNN1855, PNN1815, PNN1707);
not NOT1_548 (PNN1856, PNN1815);
not NOT1_549 (PNN1857, PNN1818);
nand NAND2_550 (PNN1858, PNN1798, PNN290);
not NOT1_551 (PNN1864, PNN1812);
nand NAND2_552 (PNN1865, PNN1812, PNN1728);
buf BUFF1_553 (PNN1866, PNN1798);
buf BUFF1_554 (PNN1869, PNN1802);
buf BUFF1_555 (PNN1872, PNN1802);
nand NAND2_556 (PNN1875, PNN1808, PNN1837);
nand NAND2_557 (PNN1878, PNN1821, PNN1848);
nand NAND2_558 (PNN1879, PNN1823, PNN1849);
nand NAND2_559 (PNN1882, PNN1841, PNN1768);
not NOT1_560 (PNN1883, PNN1841);
nand NAND2_561 (PNN1884, PNN1826, PNN1852);
nand NAND2_562 (PNN1885, PNN1643, PNN1856);
nand NAND2_563 (PNN1889, PNN1830, PNN290);
not NOT1_564 (PNN1895, PNN1838);
nand NAND2_565 (PNN1896, PNN1838, PNN1785);
nand NAND2_566 (PNN1897, PNN1640, PNN1864);
not NOT1_567 (PNN1898, PNN1850);
buf BUFF1_568 (PNN1902, PNN1830);
not NOT1_569 (PNN1910, PNN1878);
nand NAND2_570 (PNN1911, PNN1717, PNN1883);
not NOT1_571 (PNN1912, PNN1884);
nand NAND2_572 (PNN1913, PNN1855, PNN1885);
not NOT1_573 (PNN1915, PNN1866);
nand NAND2_574 (PNN1919, PNN1872, PNN919);
not NOT1_575 (PNN1920, PNN1872);
nand NAND2_576 (PNN1921, PNN1869, PNN920);
not NOT1_577 (PNN1922, PNN1869);
not NOT1_578 (PNN1923, PNN1875);
nand NAND2_579 (PNN1924, PNN1714, PNN1895);
buf BUFF1_580 (PNN1927, PNN1858);
buf BUFF1_581 (PNN1930, PNN1858);
nand NAND2_582 (PNN1933, PNN1865, PNN1897);
nand NAND2_583 (PNN1936, PNN1882, PNN1911);
not NOT1_584 (PNN1937, PNN1898);
not NOT1_585 (PNN1938, PNN1902);
nand NAND2_586 (PNN1941, PNN679, PNN1920);
nand NAND2_587 (PNN1942, PNN676, PNN1922);
buf BUFF1_588 (PNN1944, PNN1879);
not NOT1_589 (PNN1947, PNN1913);
buf BUFF1_590 (PNN1950, PNN1889);
buf BUFF1_591 (PNN1953, PNN1889);
buf BUFF1_592 (PNN1958, PNN1879);
nand NAND2_593 (PNN1961, PNN1896, PNN1924);
and AND2_594 (PNN1965, PNN1910, PNN601);
and AND2_595 (PNN1968, PNN602, PNN1912);
nand NAND2_596 (PNN1975, PNN1930, PNN917);
not NOT1_597 (PNN1976, PNN1930);
nand NAND2_598 (PNN1977, PNN1927, PNN918);
not NOT1_599 (PNN1978, PNN1927);
nand NAND2_600 (PNN1979, PNN1919, PNN1941);
nand NAND2_601 (PNN1980, PNN1921, PNN1942);
not NOT1_602 (PNN1985, PNN1933);
not NOT1_603 (PNN1987, PNN1936);
not NOT1_604 (PNN1999, PNN1944);
nand NAND2_605 (PNN2000, PNN1944, PNN1937);
not NOT1_606 (PNN2002, PNN1947);
nand NAND2_607 (PNN2003, PNN1947, PNN1499);
nand NAND2_608 (PNN2004, PNN1953, PNN1350);
not NOT1_609 (PNN2005, PNN1953);
nand NAND2_610 (PNN2006, PNN1950, PNN1351);
not NOT1_611 (PNN2007, PNN1950);
nand NAND2_612 (PNN2008, PNN673, PNN1976);
nand NAND2_613 (PNN2009, PNN670, PNN1978);
not NOT1_614 (PNN2012, PNN1979);
not NOT1_615 (PNN2013, PNN1958);
nand NAND2_616 (PNN2014, PNN1958, PNN1923);
not NOT1_617 (PNN2015, PNN1961);
nand NAND2_618 (PNN2016, PNN1961, PNN1635);
not NOT1_619 (PNN2018, PNN1965);
not NOT1_620 (PNN2019, PNN1968);
nand NAND2_621 (PNN2020, PNN1898, PNN1999);
not NOT1_622 (PNN2021, PNN1987);
nand NAND2_623 (PNN2022, PNN1987, PNN1591);
nand NAND2_624 (PNN2023, PNN1440, PNN2002);
nand NAND2_625 (PNN2024, PNN1261, PNN2005);
nand NAND2_626 (PNN2025, PNN1258, PNN2007);
nand NAND2_627 (PNN2026, PNN1975, PNN2008);
nand NAND2_628 (PNN2027, PNN1977, PNN2009);
not NOT1_629 (PNN2030, PNN1980);
buf BUFF1_630 (PNN2033, PNN1980);
nand NAND2_631 (PNN2036, PNN1875, PNN2013);
nand NAND2_632 (PNN2037, PNN1571, PNN2015);
nand NAND2_633 (PNN2038, PNN2020, PNN2000);
nand NAND2_634 (PNN2039, PNN1534, PNN2021);
nand NAND2_635 (PNN2040, PNN2023, PNN2003);
nand NAND2_636 (PNN2041, PNN2004, PNN2024);
nand NAND2_637 (PNN2042, PNN2006, PNN2025);
not NOT1_638 (PNN2047, PNN2026);
nand NAND2_639 (PNN2052, PNN2036, PNN2014);
nand NAND2_640 (PNN2055, PNN2037, PNN2016);
not NOT1_641 (PNN2060, PNN2038);
nand NAND2_642 (PNN2061, PNN2039, PNN2022);
nand NAND2_643 (PNN2062, PNN2040, PNN290);
not NOT1_644 (PNN2067, PNN2041);
not NOT1_645 (PNN2068, PNN2027);
buf BUFF1_646 (PNN2071, PNN2027);
not NOT1_647 (PNN2076, PNN2052);
not NOT1_648 (PNN2077, PNN2055);
nand NAND2_649 (PNN2078, PNN2060, PNN290);
nand NAND2_650 (PNN2081, PNN2061, PNN290);
not NOT1_651 (PNN2086, PNN2042);
buf BUFF1_652 (PNN2089, PNN2042);
and AND2_653 (PNN2104, PNN2030, PNN2068);
and AND2_654 (PNN2119, PNN2033, PNN2068);
and AND2_655 (PNN2129, PNN2030, PNN2071);
and AND2_656 (PNN2143, PNN2033, PNN2071);
buf BUFF1_657 (PNN2148, PNN2062);
buf BUFF1_658 (PNN2151, PNN2062);
buf BUFF1_659 (PNN2196, PNN2078);
buf BUFF1_660 (PNN2199, PNN2078);
buf BUFF1_661 (PNN2202, PNN2081);
buf BUFF1_662 (PNN2205, PNN2081);
nand NAND2_663 (PNN2214, PNN2151, PNN915);
not NOT1_664 (PNN2215, PNN2151);
nand NAND2_665 (PNN2216, PNN2148, PNN916);
not NOT1_666 (PNN2217, PNN2148);
nand NAND2_667 (PNN2222, PNN2199, PNN1348);
not NOT1_668 (PNN2223, PNN2199);
nand NAND2_669 (PNN2224, PNN2196, PNN1349);
not NOT1_670 (PNN2225, PNN2196);
nand NAND2_671 (PNN2226, PNN2205, PNN913);
not NOT1_672 (PNN2227, PNN2205);
nand NAND2_673 (PNN2228, PNN2202, PNN914);
not NOT1_674 (PNN2229, PNN2202);
nand NAND2_675 (PNN2230, PNN667, PNN2215);
nand NAND2_676 (PNN2231, PNN664, PNN2217);
nand NAND2_677 (PNN2232, PNN1255, PNN2223);
nand NAND2_678 (PNN2233, PNN1252, PNN2225);
nand NAND2_679 (PNN2234, PNN661, PNN2227);
nand NAND2_680 (PNN2235, PNN658, PNN2229);
nand NAND2_681 (PNN2236, PNN2214, PNN2230);
nand NAND2_682 (PNN2237, PNN2216, PNN2231);
nand NAND2_683 (PNN2240, PNN2222, PNN2232);
nand NAND2_684 (PNN2241, PNN2224, PNN2233);
nand NAND2_685 (PNN2244, PNN2226, PNN2234);
nand NAND2_686 (PNN2245, PNN2228, PNN2235);
not NOT1_687 (PNN2250, PNN2236);
not NOT1_688 (PNN2253, PNN2240);
not NOT1_689 (PNN2256, PNN2244);
not NOT1_690 (PNN2257, PNN2237);
buf BUFF1_691 (PNN2260, PNN2237);
not NOT1_692 (PNN2263, PNN2241);
and AND2_693 (PNN2266, PNN1164, PNN2241);
not NOT1_694 (PNN2269, PNN2245);
and AND2_695 (PNN2272, PNN1168, PNN2245);
nand NAND8_696 (PNN2279, PNN2067, PNN2012, PNN2047, PNN2250, PNN899, PNN2256, PNN2253, PNN903);
buf BUFF1_697 (PNN2286, PNN2266);
buf BUFF1_698 (PNN2297, PNN2266);
buf BUFF1_699 (PNN2315, PNN2272);
buf BUFF1_700 (PNN2326, PNN2272);
and AND2_701 (PNN2340, PNN2086, PNN2257);
and AND2_702 (PNN2353, PNN2089, PNN2257);
and AND2_703 (PNN2361, PNN2086, PNN2260);
and AND2_704 (PNN2375, PNN2089, PNN2260);
and AND4_705 (PNN2384, PNN338, PNN2279, PNN313, PNN313);
and AND2_706 (PNN2385, PNN1163, PNN2263);
and AND2_707 (PNN2386, PNN1164, PNN2263);
and AND2_708 (PNN2426, PNN1167, PNN2269);
and AND2_709 (PNN2427, PNN1168, PNN2269);
nand NAND5_710 (PNN2537, PNN2286, PNN2315, PNN2361, PNN2104, PNN1171);
nand NAND5_711 (PNN2540, PNN2286, PNN2315, PNN2340, PNN2129, PNN1171);
nand NAND5_712 (PNN2543, PNN2286, PNN2315, PNN2340, PNN2119, PNN1171);
nand NAND5_713 (PNN2546, PNN2286, PNN2315, PNN2353, PNN2104, PNN1171);
nand NAND5_714 (PNN2549, PNN2297, PNN2315, PNN2375, PNN2119, PNN1188);
nand NAND5_715 (PNN2552, PNN2297, PNN2326, PNN2361, PNN2143, PNN1188);
nand NAND5_716 (PNN2555, PNN2297, PNN2326, PNN2375, PNN2129, PNN1188);
and AND5_717 (PNN2558, PNN2286, PNN2315, PNN2361, PNN2104, PNN1171);
and AND5_718 (PNN2561, PNN2286, PNN2315, PNN2340, PNN2129, PNN1171);
and AND5_719 (PNN2564, PNN2286, PNN2315, PNN2340, PNN2119, PNN1171);
and AND5_720 (PNN2567, PNN2286, PNN2315, PNN2353, PNN2104, PNN1171);
and AND5_721 (PNN2570, PNN2297, PNN2315, PNN2375, PNN2119, PNN1188);
and AND5_722 (PNN2573, PNN2297, PNN2326, PNN2361, PNN2143, PNN1188);
and AND5_723 (PNN2576, PNN2297, PNN2326, PNN2375, PNN2129, PNN1188);
nand NAND5_724 (PNN2594, PNN2286, PNN2427, PNN2361, PNN2129, PNN1171);
nand NAND5_725 (PNN2597, PNN2297, PNN2427, PNN2361, PNN2119, PNN1171);
nand NAND5_726 (PNN2600, PNN2297, PNN2427, PNN2375, PNN2104, PNN1171);
nand NAND5_727 (PNN2603, PNN2297, PNN2427, PNN2340, PNN2143, PNN1171);
nand NAND5_728 (PNN2606, PNN2297, PNN2427, PNN2353, PNN2129, PNN1188);
nand NAND5_729 (PNN2611, PNN2386, PNN2326, PNN2361, PNN2129, PNN1188);
nand NAND5_730 (PNN2614, PNN2386, PNN2326, PNN2361, PNN2119, PNN1188);
nand NAND5_731 (PNN2617, PNN2386, PNN2326, PNN2375, PNN2104, PNN1188);
nand NAND5_732 (PNN2620, PNN2386, PNN2326, PNN2353, PNN2129, PNN1188);
nand NAND5_733 (PNN2627, PNN2297, PNN2427, PNN2340, PNN2104, PNN926);
nand NAND5_734 (PNN2628, PNN2386, PNN2326, PNN2340, PNN2104, PNN926);
nand NAND5_735 (PNN2629, PNN2386, PNN2427, PNN2361, PNN2104, PNN926);
nand NAND5_736 (PNN2630, PNN2386, PNN2427, PNN2340, PNN2129, PNN926);
nand NAND5_737 (PNN2631, PNN2386, PNN2427, PNN2340, PNN2119, PNN926);
nand NAND5_738 (PNN2632, PNN2386, PNN2427, PNN2353, PNN2104, PNN926);
nand NAND5_739 (PNN2633, PNN2386, PNN2426, PNN2340, PNN2104, PNN926);
nand NAND5_740 (PNN2634, PNN2385, PNN2427, PNN2340, PNN2104, PNN926);
and AND5_741 (PNN2639, PNN2286, PNN2427, PNN2361, PNN2129, PNN1171);
and AND5_742 (PNN2642, PNN2297, PNN2427, PNN2361, PNN2119, PNN1171);
and AND5_743 (PNN2645, PNN2297, PNN2427, PNN2375, PNN2104, PNN1171);
and AND5_744 (PNN2648, PNN2297, PNN2427, PNN2340, PNN2143, PNN1171);
and AND5_745 (PNN2651, PNN2297, PNN2427, PNN2353, PNN2129, PNN1188);
and AND5_746 (PNN2655, PNN2386, PNN2326, PNN2361, PNN2129, PNN1188);
and AND5_747 (PNN2658, PNN2386, PNN2326, PNN2361, PNN2119, PNN1188);
and AND5_748 (PNN2661, PNN2386, PNN2326, PNN2375, PNN2104, PNN1188);
and AND5_749 (PNN2664, PNN2386, PNN2326, PNN2353, PNN2129, PNN1188);
nand NAND2_750 (PNN2669, PNN2558, PNN534);
not NOT1_751 (PNN2670, PNN2558);
nand NAND2_752 (PNN2671, PNN2561, PNN535);
not NOT1_753 (PNN2672, PNN2561);
nand NAND2_754 (PNN2673, PNN2564, PNN536);
not NOT1_755 (PNN2674, PNN2564);
nand NAND2_756 (PNN2675, PNN2567, PNN537);
not NOT1_757 (PNN2676, PNN2567);
nand NAND2_758 (PNN2682, PNN2570, PNN543);
not NOT1_759 (PNN2683, PNN2570);
nand NAND2_760 (PNN2688, PNN2573, PNN548);
not NOT1_761 (PNN2689, PNN2573);
nand NAND2_762 (PNN2690, PNN2576, PNN549);
not NOT1_763 (PNN2691, PNN2576);
and AND8_764 (PNN2710, PNN2627, PNN2628, PNN2629, PNN2630, PNN2631, PNN2632, PNN2633, PNN2634);
nand NAND2_765 (PNN2720, PNN343, PNN2670);
nand NAND2_766 (PNN2721, PNN346, PNN2672);
nand NAND2_767 (PNN2722, PNN349, PNN2674);
nand NAND2_768 (PNN2723, PNN352, PNN2676);
nand NAND2_769 (PNN2724, PNN2639, PNN538);
not NOT1_770 (PNN2725, PNN2639);
nand NAND2_771 (PNN2726, PNN2642, PNN539);
not NOT1_772 (PNN2727, PNN2642);
nand NAND2_773 (PNN2728, PNN2645, PNN540);
not NOT1_774 (PNN2729, PNN2645);
nand NAND2_775 (PNN2730, PNN2648, PNN541);
not NOT1_776 (PNN2731, PNN2648);
nand NAND2_777 (PNN2732, PNN2651, PNN542);
not NOT1_778 (PNN2733, PNN2651);
nand NAND2_779 (PNN2734, PNN370, PNN2683);
nand NAND2_780 (PNN2735, PNN2655, PNN544);
not NOT1_781 (PNN2736, PNN2655);
nand NAND2_782 (PNN2737, PNN2658, PNN545);
not NOT1_783 (PNN2738, PNN2658);
nand NAND2_784 (PNN2739, PNN2661, PNN546);
not NOT1_785 (PNN2740, PNN2661);
nand NAND2_786 (PNN2741, PNN2664, PNN547);
not NOT1_787 (PNN2742, PNN2664);
nand NAND2_788 (PNN2743, PNN385, PNN2689);
nand NAND2_789 (PNN2744, PNN388, PNN2691);
nand NAND8_790 (PNN2745, PNN2537, PNN2540, PNN2543, PNN2546, PNN2594, PNN2597, PNN2600, PNN2603);
nand NAND8_791 (PNN2746, PNN2606, PNN2549, PNN2611, PNN2614, PNN2617, PNN2620, PNN2552, PNN2555);
and AND8_792 (PNN2747, PNN2537, PNN2540, PNN2543, PNN2546, PNN2594, PNN2597, PNN2600, PNN2603);
and AND8_793 (PNN2750, PNN2606, PNN2549, PNN2611, PNN2614, PNN2617, PNN2620, PNN2552, PNN2555);
nand NAND2_794 (PNN2753, PNN2669, PNN2720);
nand NAND2_795 (PNN2754, PNN2671, PNN2721);
nand NAND2_796 (PNN2755, PNN2673, PNN2722);
nand NAND2_797 (PNN2756, PNN2675, PNN2723);
nand NAND2_798 (PNN2757, PNN355, PNN2725);
nand NAND2_799 (PNN2758, PNN358, PNN2727);
nand NAND2_800 (PNN2759, PNN361, PNN2729);
nand NAND2_801 (PNN2760, PNN364, PNN2731);
nand NAND2_802 (PNN2761, PNN367, PNN2733);
nand NAND2_803 (PNN2762, PNN2682, PNN2734);
nand NAND2_804 (PNN2763, PNN373, PNN2736);
nand NAND2_805 (PNN2764, PNN376, PNN2738);
nand NAND2_806 (PNN2765, PNN379, PNN2740);
nand NAND2_807 (PNN2766, PNN382, PNN2742);
nand NAND2_808 (PNN2767, PNN2688, PNN2743);
nand NAND2_809 (PNN2768, PNN2690, PNN2744);
and AND2_810 (PNN2773, PNN2745, PNN275);
and AND2_811 (PNN2776, PNN2746, PNN276);
nand NAND2_812 (PNN2779, PNN2724, PNN2757);
nand NAND2_813 (PNN2780, PNN2726, PNN2758);
nand NAND2_814 (PNN2781, PNN2728, PNN2759);
nand NAND2_815 (PNN2782, PNN2730, PNN2760);
nand NAND2_816 (PNN2783, PNN2732, PNN2761);
nand NAND2_817 (PNN2784, PNN2735, PNN2763);
nand NAND2_818 (PNN2785, PNN2737, PNN2764);
nand NAND2_819 (PNN2786, PNN2739, PNN2765);
nand NAND2_820 (PNN2787, PNN2741, PNN2766);
and AND3_821 (PNN2788, PNN2747, PNN2750, PNN2710);
nand NAND2_822 (PNN2789, PNN2747, PNN2750);
and AND4_823 (PNN2800, PNN338, PNN2279, PNN99, PNN2788);
nand NAND2_824 (PNN2807, PNN2773, PNN2018);
not NOT1_825 (PNN2808, PNN2773);
nand NAND2_826 (PNN2809, PNN2776, PNN2019);
not NOT1_827 (PNN2810, PNN2776);
nor NOR2_828 (PNN2811, PNN2384, PNN2800);
and AND3_829 (PNN2812, PNN897, PNN283, PNN2789);
and AND3_830 (PNN2815, PNN76, PNN283, PNN2789);
and AND3_831 (PNN2818, PNN82, PNN283, PNN2789);
and AND3_832 (PNN2821, PNN85, PNN283, PNN2789);
and AND3_833 (PNN2824, PNN898, PNN283, PNN2789);
nand NAND2_834 (PNN2827, PNN1965, PNN2808);
nand NAND2_835 (PNN2828, PNN1968, PNN2810);
and AND3_836 (PNN2829, PNN79, PNN283, PNN2789);
nand NAND2_837 (PNN2843, PNN2807, PNN2827);
nand NAND2_838 (PNN2846, PNN2809, PNN2828);
nand NAND2_839 (PNN2850, PNN2812, PNN2076);
nand NAND2_840 (PNN2851, PNN2815, PNN2077);
nand NAND2_841 (PNN2852, PNN2818, PNN1915);
nand NAND2_842 (PNN2853, PNN2821, PNN1857);
nand NAND2_843 (PNN2854, PNN2824, PNN1938);
not NOT1_844 (PNN2857, PNN2812);
not NOT1_845 (PNN2858, PNN2815);
not NOT1_846 (PNN2859, PNN2818);
not NOT1_847 (PNN2860, PNN2821);
not NOT1_848 (PNN2861, PNN2824);
not NOT1_849 (PNN2862, PNN2829);
nand NAND2_850 (PNN2863, PNN2829, PNN1985);
nand NAND2_851 (PNN2866, PNN2052, PNN2857);
nand NAND2_852 (PNN2867, PNN2055, PNN2858);
nand NAND2_853 (PNN2868, PNN1866, PNN2859);
nand NAND2_854 (PNN2869, PNN1818, PNN2860);
nand NAND2_855 (PNN2870, PNN1902, PNN2861);
nand NAND2_856 (PNN2871, PNN2843, PNN886);
not NOT1_857 (PNN2872, PNN2843);
nand NAND2_858 (PNN2873, PNN2846, PNN887);
not NOT1_859 (PNN2874, PNN2846);
nand NAND2_860 (PNN2875, PNN1933, PNN2862);
nand NAND2_861 (PNN2876, PNN2866, PNN2850);
nand NAND2_862 (PNN2877, PNN2867, PNN2851);
nand NAND2_863 (PNN2878, PNN2868, PNN2852);
nand NAND2_864 (PNN2879, PNN2869, PNN2853);
nand NAND2_865 (PNN2880, PNN2870, PNN2854);
nand NAND2_866 (PNN2881, PNN682, PNN2872);
nand NAND2_867 (PNN2882, PNN685, PNN2874);
nand NAND2_868 (PNN2883, PNN2875, PNN2863);
and AND2_869 (PNN2886, PNN2876, PNN550);
and AND2_870 (PNN2887, PNN551, PNN2877);
and AND2_871 (PNN2888, PNN553, PNN2878);
and AND2_872 (PNN2889, PNN2879, PNN554);
and AND2_873 (PNN2890, PNN555, PNN2880);
nand NAND2_874 (PNN2891, PNN2871, PNN2881);
nand NAND2_875 (PNN2892, PNN2873, PNN2882);
nand NAND2_876 (PNN2895, PNN2883, PNN1461);
not NOT1_877 (PNN2896, PNN2883);
nand NAND2_878 (PNN2897, PNN1383, PNN2896);
nand NAND2_879 (PNN2898, PNN2895, PNN2897);
and AND2_880 (PNN2899, PNN2898, PNN552);

endmodule


module c1908_clk_ipFF (clk,PNN1,PNN4,PNN7,PNN10,PNN13,PNN16,PNN19,PNN22,PNN25,PNN28,
              PNN31,PNN34,PNN37,PNN40,PNN43,PNN46,PNN49,PNN53,PNN56,PNN60,
              PNN63,PNN66,PNN69,PNN72,PNN76,PNN79,PNN82,PNN85,PNN88,PNN91,
              PNN94,PNN99,PNN104,Q_PNN2753,Q_PNN2754,Q_PNN2755,Q_PNN2756,Q_PNN2762,Q_PNN2767,Q_PNN2768,
              Q_PNN2779,Q_PNN2780,Q_PNN2781,Q_PNN2782,Q_PNN2783,Q_PNN2784,Q_PNN2785,Q_PNN2786,Q_PNN2787,Q_PNN2811,
              Q_PNN2886,Q_PNN2887,Q_PNN2888,Q_PNN2889,Q_PNN2890,Q_PNN2891,Q_PNN2892,Q_PNN2899);

input clk,PNN1,PNN4,PNN7,PNN10,PNN13,PNN16,PNN19,PNN22,PNN25,PNN28,
      PNN31,PNN34,PNN37,PNN40,PNN43,PNN46,PNN49,PNN53,PNN56,PNN60,
      PNN63,PNN66,PNN69,PNN72,PNN76,PNN79,PNN82,PNN85,PNN88,PNN91,
      PNN94,PNN99,PNN104;

output Q_PNN2753,Q_PNN2754,Q_PNN2755,Q_PNN2756,Q_PNN2762,Q_PNN2767,Q_PNN2768,Q_PNN2779,Q_PNN2780,Q_PNN2781,
       Q_PNN2782,Q_PNN2783,Q_PNN2784,Q_PNN2785,Q_PNN2786,Q_PNN2787,Q_PNN2811,Q_PNN2886,Q_PNN2887,Q_PNN2888,
       Q_PNN2889,Q_PNN2890,Q_PNN2891,Q_PNN2892,Q_PNN2899;


 c1908 C_0(IN_PNN1,IN_PNN4,IN_PNN7,IN_PNN10,IN_PNN13,IN_PNN16,IN_PNN19,IN_PNN22,IN_PNN25,IN_PNN28,
              IN_PNN31,IN_PNN34,IN_PNN37,IN_PNN40,IN_PNN43,IN_PNN46,IN_PNN49,IN_PNN53,IN_PNN56,IN_PNN60,
              IN_PNN63,IN_PNN66,IN_PNN69,IN_PNN72,IN_PNN76,IN_PNN79,IN_PNN82,IN_PNN85,IN_PNN88,IN_PNN91,
              IN_PNN94,IN_PNN99,IN_PNN104,PNN2753,PNN2754,PNN2755,PNN2756,PNN2762,PNN2767,PNN2768,
              PNN2779,PNN2780,PNN2781,PNN2782,PNN2783,PNN2784,PNN2785,PNN2786,PNN2787,PNN2811,
              PNN2886,PNN2887,PNN2888,PNN2889,PNN2890,PNN2891,PNN2892,PNN2899);



//input FFs
dff iDFF_1 (IN_PNN1,  PNN1, clk);
dff iDFF_2 (IN_PNN4,  PNN4, clk);
dff iDFF_3 (IN_PNN7,  PNN7, clk);
dff iDFF_4 (IN_PNN10, PNN10, clk);
dff iDFF_5 (IN_PNN13, PNN13, clk);
dff iDFF_6 (IN_PNN16, PNN16, clk);
dff iDFF_7 (IN_PNN19, PNN19, clk);
dff iDFF_8 (IN_PNN22, PNN22, clk);
dff iDFF_9 (IN_PNN25, PNN25, clk);
dff iDFF_10(IN_PNN28, PNN28, clk);
dff iDFF_11(IN_PNN31, PNN31, clk);
dff iDFF_12(IN_PNN34, PNN34, clk);
dff iDFF_13(IN_PNN37, PNN37, clk);
dff iDFF_14(IN_PNN40, PNN40, clk);
dff iDFF_15(IN_PNN43, PNN43, clk);
dff iDFF_16(IN_PNN46, PNN46, clk);
dff iDFF_17(IN_PNN49, PNN49, clk);
dff iDFF_18(IN_PNN53, PNN53, clk);
dff iDFF_19(IN_PNN56, PNN56, clk);
dff iDFF_20(IN_PNN60, PNN60, clk);
dff iDFF_21(IN_PNN63, PNN63, clk);
dff iDFF_22(IN_PNN66, PNN66, clk);
dff iDFF_23(IN_PNN69, PNN69, clk);
dff iDFF_24(IN_PNN72, PNN72, clk);
dff iDFF_25(IN_PNN76, PNN76, clk);
dff iDFF_26(IN_PNN79, PNN79, clk);
dff iDFF_27(IN_PNN82, PNN82, clk);
dff iDFF_28(IN_PNN85, PNN85, clk);
dff iDFF_29(IN_PNN88, PNN88, clk);
dff iDFF_30(IN_PNN91, PNN91, clk);
dff iDFF_31(IN_PNN94, PNN94, clk);
dff iDFF_32(IN_PNN99, PNN99, clk);
dff iDFF_33(IN_PNN104, PNN104,clk);


//output FFs	
  dff DFF_0(Q_PNN2753,PNN2753,clk);
  dff DFF_1(Q_PNN2754,PNN2754,clk);
  dff DFF_2(Q_PNN2755,PNN2755,clk);
  dff DFF_3(Q_PNN2756,PNN2756,clk);
  dff DFF_4(Q_PNN2762,PNN2762,clk);
  dff DFF_5(Q_PNN2767,PNN2767,clk);
  dff DFF_6(Q_PNN2768,PNN2768,clk);
  dff DFF_7(Q_PNN2779,PNN2779,clk);
  dff DFF_8(Q_PNN2780,PNN2780,clk);
  dff DFF_9(Q_PNN2781,PNN2781,clk);
  dff DFF_10(Q_PNN2782,PNN2782,clk);
  dff DFF_11(Q_PNN2783,PNN2783,clk);
  dff DFF_12(Q_PNN2784,PNN2784,clk);
  dff DFF_13(Q_PNN2785,PNN2785,clk);
  dff DFF_14(Q_PNN2786,PNN2786,clk);
  dff DFF_15(Q_PNN2787,PNN2787,clk);
  dff DFF_16(Q_PNN2811,PNN2811,clk);
  dff DFF_17(Q_PNN2886,PNN2886,clk);
  dff DFF_18(Q_PNN2887,PNN2887,clk);
  dff DFF_19(Q_PNN2888,PNN2888,clk);
  dff DFF_20(Q_PNN2889,PNN2889,clk);
  dff DFF_21(Q_PNN2890,PNN2890,clk);
  dff DFF_22(Q_PNN2891,PNN2891,clk);
  dff DFF_23(Q_PNN2892,PNN2892,clk);
  dff DFF_24(Q_PNN2899,PNN2899,clk);


endmodule



