**clk_4227_glitch_1.66344711153e-09_random_gate_HS65_GS_DFPQX9_random_drain_21_deck_number_1
****Template spice file***

.include  ../hspice_glitch_CORE65GPSVT_selected_lib_vg.sp
.include /home/users/nanditha/Documents/utility/65nm/hspice_65nm_models/diodeiso_typ.txt
.include /home/users/nanditha/Documents/utility/65nm/hspice_65nm_models/ptm_nmos_65_no_X.txt
.include /home/users/nanditha/Documents/utility/65nm/hspice_65nm_models/ptm_pmos_65_no_X.txt
**********Subckt begins*********

.SUBCKT c499_clk_opFF 
+ clk PNN1 PNN5 PNN9 PNN13 PNN17 PNN21 PNN25 PNN29 PNN33 
+ PNN37 PNN41 PNN45 PNN49 PNN53 PNN57 PNN61 PNN65 PNN69 PNN73 
+ PNN77 PNN81 PNN85 PNN89 PNN93 PNN97 PNN101 PNN105 PNN109 PNN113 
+ PNN117 PNN121 PNN125 PNN129 PNN130 PNN131 PNN132 PNN133 PNN134 PNN135 
+ PNN136 PNN137 Qout_PNN724 Qout_PNN725 Qout_PNN726 Qout_PNN727 Qout_PNN728 Qout_PNN729 Qout_PNN730 Qout_PNN731 
+ Qout_PNN732 Qout_PNN733 Qout_PNN734 Qout_PNN735 Qout_PNN736 Qout_PNN737 Qout_PNN738 Qout_PNN739 Qout_PNN740 Qout_PNN741 
+ Qout_PNN742 Qout_PNN743 Qout_PNN744 Qout_PNN745 Qout_PNN746 Qout_PNN747 Qout_PNN748 Qout_PNN749 Qout_PNN750 Qout_PNN751 
+ Qout_PNN752 Qout_PNN753 Qout_PNN754 Qout_PNN755 

C1_255 U298:A 0 0.000031PF
C2_255 clk_r_REG32_S2:Q 0 0.000031PF
R1_255 U298:A clk_r_REG32_S2:Q 0.304000

C1_183 U228:Z 0 0.000111PF
C2_183 U258:A 0 0.000111PF
R1_183 U258:A U228:Z 0.912000

C1_241 U270:A 0 0.000107PF
C2_241 clk_r_REG46_S2:Q 0 0.000107PF
R1_241 U270:A clk_r_REG46_S2:Q 1.064000

C1_222 clk_r_REG50_S2:Q 0 0.000399PF
C2_222 U262:A 0 0.000399PF
R1_222 U262:A clk_r_REG50_S2:Q 3.496000

C1_212 U260:A 0 0.000076PF
C2_212 clk_r_REG51_S2:Q 0 0.000076PF
R1_212 U260:A clk_r_REG51_S2:Q 0.760000

C1_265 clk_r_REG21_S2:Q 0 0.000045PF
C2_265 n43_4 0 0.000141PF
C3_265 n43_3 0 0.000141PF
C4_265 n43_2 0 0.000201PF
C5_265 U313:A 0 0.000178PF
R1_265 n43_2 U313:A 1.976000
R2_265 n43_2 n43_3 4.000000
R3_265 n43_4 n43_3 1.520000
R4_265 n43_4 clk_r_REG21_S2:Q 4.000000

C1_268 clk_r_REG7_S2:Q 0 0.000045PF
C2_268 n46_4 0 0.000148PF
C3_268 n46_3 0 0.000148PF
C4_268 n46_2 0 0.000105PF
C5_268 oDFF_8_q_reg:D 0 0.000082PF
R1_268 n46_2 oDFF_8_q_reg:D 0.912000
R2_268 n46_2 n46_3 4.000000
R3_268 n46_3 n46_4 1.672000
R4_268 n46_4 clk_r_REG7_S2:Q 4.000000

C1_111 oDFF_29_q_reg:D 0 0.000045PF
C2_111 Q_PNN752_3 0 0.000090PF
C3_111 Q_PNN752_2 0 0.000090PF
C4_111 U266:Z 0 0.000045PF
R1_111 U266:Z Q_PNN752_2 4.000000
R2_111 Q_PNN752_2 Q_PNN752_3 1.520000
R3_111 Q_PNN752_3 oDFF_29_q_reg:D 4.000000

C1_264 clk_r_REG22_S2:Q 0 0.000045PF
C2_264 n42_4 0 0.000146PF
C3_264 n42_3 0 0.000146PF
C4_264 n42_2 0 0.000290PF
C5_264 U314:A 0 0.000268PF
R1_264 n42_2 U314:A 2.888000
R2_264 n42_2 n42_3 4.000000
R3_264 n42_4 n42_3 1.520000
R4_264 n42_4 clk_r_REG22_S2:Q 4.000000

C1_86 clk_r_REG8_S2:D 0 0.000045PF
C2_86 Q_PNN727_5 0 0.000068PF
C3_86 Q_PNN727_4 0 0.000102PF
C4_86 Q_PNN727_3 0 0.000110PF
C5_86 Q_PNN727_2 0 0.000076PF
C6_86 U240:Z 0 0.000045PF
R1_86 U240:Z Q_PNN727_2 4.000000
R2_86 Q_PNN727_2 Q_PNN727_3 0.912000
R3_86 Q_PNN727_3 Q_PNN727_4 0.152000
R4_86 Q_PNN727_4 Q_PNN727_5 1.064000
R5_86 Q_PNN727_5 clk_r_REG8_S2:D 4.000000

C1_107 U274:Z 0 0.000045PF
C2_107 Q_PNN748_4 0 0.000082PF
C3_107 Q_PNN748_3 0 0.000082PF
C4_107 Q_PNN748_2 0 0.000122PF
C5_107 oDFF_25_q_reg:D 0 0.000099PF
R1_107 oDFF_25_q_reg:D Q_PNN748_2 1.064000
R2_107 Q_PNN748_2 Q_PNN748_3 4.000000
R3_107 Q_PNN748_4 Q_PNN748_3 1.368000
R4_107 Q_PNN748_4 U274:Z 4.000000

C1_308 U275:Z 0 0.000045PF
C2_308 n82_3 0 0.000187PF
C3_308 n82_2 0 0.000187PF
C4_308 U274:B 0 0.000045PF
R1_308 U274:B n82_2 4.000000
R2_308 n82_3 n82_2 1.824000
R3_308 n82_3 U275:Z 4.000000

C1_151 clk_r_REG22_S2:D 0 0.000045PF
C2_151 c0_n29_4 0 0.000107PF
C3_151 c0_n29_3 0 0.000107PF
C4_151 c0_n29_2 0 0.000153PF
C5_151 U165:Z 0 0.000130PF
R1_151 c0_n29_2 U165:Z 1.064000
R2_151 c0_n29_2 c0_n29_3 4.000000
R3_151 c0_n29_3 c0_n29_4 1.368000
R4_151 c0_n29_4 clk_r_REG22_S2:D 4.000000

C1_145 oDFF_31_q_reg:Q 0 0.000045PF
C2_145 Qout_PNN754_5 0 0.002591PF
C3_145 Qout_PNN754_4 0 0.002591PF
C4_145 Qout_PNN754_3 0 0.000046PF
C5_145 Qout_PNN754_2 0 0.000046PF
C6_145 Qout_PNN754 0 0.000042PF
R1_145 Qout_PNN754 Qout_PNN754_2 4.000000
R2_145 Qout_PNN754_3 Qout_PNN754_2 0.304000
R3_145 Qout_PNN754_3 Qout_PNN754_4 4.000000
R4_145 Qout_PNN754_5 Qout_PNN754_4 32.679999
R5_145 Qout_PNN754_5 oDFF_31_q_reg:Q 4.000000

C1_307 U273:Z 0 0.000045PF
C2_307 n81_5 0 0.000169PF
C3_307 n81_4 0 0.000203PF
C4_307 n81_3 0 0.000165PF
C5_307 n81_2 0 0.000130PF
C6_307 U272:B 0 0.000045PF
R1_307 U272:B n81_2 4.000000
R2_307 n81_3 n81_2 0.912000
R3_307 n81_4 n81_3 0.152000
R4_307 n81_5 n81_4 0.912000
R5_307 n81_5 U273:Z 4.000000

C1_167 U235:Z 0 0.000045PF
C2_167 n103_3 0 0.000122PF
C3_167 n103_2 0 0.000122PF
C4_167 U234:B 0 0.000045PF
R1_167 U234:B n103_2 4.000000
R2_167 n103_2 n103_3 1.520000
R3_167 n103_3 U235:Z 4.000000

C1_263 clk_r_REG3_S2:Q 0 0.000045PF
C2_263 n41_4 0 0.000461PF
C3_263 n41_3 0 0.000461PF
C4_263 n41_2 0 0.000099PF
C5_263 U308:A 0 0.000077PF
R1_263 n41_2 U308:A 0.760000
R2_263 n41_2 n41_3 4.000000
R3_263 n41_4 n41_3 3.344000
R4_263 n41_4 clk_r_REG3_S2:Q 4.000000

C1_146 oDFF_32_q_reg:Q 0 0.000045PF
C2_146 Qout_PNN755_5 0 0.002543PF
C3_146 Qout_PNN755_4 0 0.002543PF
C4_146 Qout_PNN755_3 0 0.000046PF
C5_146 Qout_PNN755_2 0 0.000046PF
C6_146 Qout_PNN755 0 0.000042PF
R1_146 Qout_PNN755 Qout_PNN755_2 4.000000
R2_146 Qout_PNN755_3 Qout_PNN755_2 0.304000
R3_146 Qout_PNN755_3 Qout_PNN755_4 4.000000
R4_146 Qout_PNN755_5 Qout_PNN755_4 30.703999
R5_146 Qout_PNN755_5 oDFF_32_q_reg:Q 4.000000

C1_60 PNN17 0 0.003783PF
C2_60 PNN17_2 0 0.003804PF
C3_60 iDFF_5_q_reg:D 0 0.000045PF
R1_60 iDFF_5_q_reg:D PNN17_2 4.000000
R2_60 PNN17 PNN17_2 32.983999

C1_123 oDFF_9_q_reg:Q 0 0.000045PF
C2_123 Qout_PNN732_4 0 0.000327PF
C3_123 Qout_PNN732_3 0 0.000361PF
C4_123 Qout_PNN732_2 0 0.005010PF
C5_123 Qout_PNN732 0 0.004955PF
R1_123 Qout_PNN732 Qout_PNN732_2 33.287999
R2_123 Qout_PNN732_3 Qout_PNN732_2 0.152000
R3_123 Qout_PNN732_3 Qout_PNN732_4 3.344000
R4_123 Qout_PNN732_4 oDFF_9_q_reg:Q 4.000000

C1_119 oDFF_5_q_reg:Q 0 0.000045PF
C2_119 Qout_PNN728_5 0 0.003885PF
C3_119 Qout_PNN728_4 0 0.003885PF
C4_119 Qout_PNN728_3 0 0.000046PF
C5_119 Qout_PNN728_2 0 0.000046PF
C6_119 Qout_PNN728 0 0.000042PF
R1_119 Qout_PNN728 Qout_PNN728_2 4.000000
R2_119 Qout_PNN728_3 Qout_PNN728_2 0.304000
R3_119 Qout_PNN728_3 Qout_PNN728_4 4.000000
R4_119 Qout_PNN728_4 Qout_PNN728_5 30.703999
R5_119 Qout_PNN728_5 oDFF_5_q_reg:Q 4.000000

C1_178 U246:B 0 0.000045PF
C2_178 n113_3 0 0.000360PF
C3_178 n113_2 0 0.000360PF
C4_178 U247:Z 0 0.000045PF
R1_178 U247:Z n113_2 4.000000
R2_178 n113_3 n113_2 1.520000
R3_178 n113_3 U246:B 4.000000

C1_298 U261:Z 0 0.000045PF
C2_298 n73_7 0 0.000170PF
C3_298 n73_6 0 0.000170PF
C4_298 n73_5 0 0.000174PF
C5_298 n73_4 0 0.000174PF
C6_298 n73_3 0 0.000151PF
C7_298 n73_2 0 0.000151PF
C8_298 U260:B 0 0.000045PF
R1_298 U260:B n73_2 4.000000
R2_298 n73_3 n73_2 1.976000
R3_298 n73_3 n73_4 4.000000
R4_298 n73_5 n73_4 1.216000
R5_298 n73_5 n73_6 4.000000
R6_298 n73_7 n73_6 1.976000
R7_298 n73_7 U261:Z 4.000000

C1_114 U260:Z 0 0.000045PF
C2_114 Q_PNN755_4 0 0.000175PF
C3_114 Q_PNN755_3 0 0.000175PF
C4_114 Q_PNN755_2 0 0.000064PF
C5_114 oDFF_32_q_reg:D 0 0.000041PF
R1_114 oDFF_32_q_reg:D Q_PNN755_2 0.456000
R2_114 Q_PNN755_2 Q_PNN755_3 4.000000
R3_114 Q_PNN755_4 Q_PNN755_3 1.824000
R4_114 Q_PNN755_4 U260:Z 4.000000

C1_324 U299:Z 0 0.000045PF
C2_324 n97_3 0 0.000148PF
C3_324 n97_2 0 0.000148PF
C4_324 U298:B 0 0.000045PF
R1_324 U298:B n97_2 4.000000
R2_324 n97_2 n97_3 1.520000
R3_324 n97_3 U299:Z 4.000000

C1_172 U162:Z 0 0.000045PF
C2_172 n108_5 0 0.000340PF
C3_172 n108_4 0 0.000340PF
C4_172 n108_3 0 0.000082PF
C5_172 U163:B 0 0.000132PF
C6_172 U161:B 0 0.000072PF
R1_172 U161:B U163:B 0.760000
R2_172 n108_3 U163:B 0.456000
R3_172 n108_3 n108_4 4.000000
R4_172 n108_4 n108_5 1.368000
R5_172 n108_5 U162:Z 4.000000

C1_226 U239:Z 0 0.000045PF
C2_226 n163_4 0 0.000305PF
C3_226 n163_3 0 0.000305PF
C4_226 n163_2 0 0.000091PF
C5_226 U237:A 0 0.000069PF
R1_226 n163_2 U237:A 0.760000
R2_226 n163_2 n163_3 4.000000
R3_226 n163_4 n163_3 1.672000
R4_226 n163_4 U239:Z 4.000000

C1_225 U237:Z 0 0.000045PF
C2_225 n162_6 0 0.000529PF
C3_225 n162_5 0 0.000564PF
C4_225 n162_4 0 0.000249PF
C5_225 n162_3 0 0.000249PF
C6_225 n162_2 0 0.000086PF
C7_225 U236:C 0 0.000045PF
R1_225 U236:C n162_2 4.000000
R2_225 n162_3 n162_2 0.152000
R3_225 n162_4 n162_3 1.976000
R4_225 n162_5 n162_4 0.152000
R5_225 n162_6 n162_5 3.648000
R6_225 n162_6 U237:Z 4.000000

C1_296 U166:D 0 0.000045PF
C2_296 n71_4 0 0.000092PF
C3_296 n71_3 0 0.000092PF
C4_296 n71_2 0 0.000060PF
C5_296 U167:Z 0 0.000037PF
R1_296 n71_2 U167:Z 0.304000
R2_296 n71_2 n71_3 4.000000
R3_296 n71_4 n71_3 1.520000
R4_296 n71_4 U166:D 4.000000

C1_260 clk_r_REG18_S2:Q 0 0.000045PF
C2_260 n39_3 0 0.000201PF
C3_260 n39_2 0 0.000201PF
C4_260 U211:A 0 0.000045PF
R1_260 U211:A n39_2 4.000000
R2_260 n39_2 n39_3 1.520000
R3_260 n39_3 clk_r_REG18_S2:Q 4.000000

C1_64 PNN33 0 0.003011PF
C2_64 PNN33_2 0 0.003032PF
C3_64 iDFF_9_q_reg:D 0 0.000045PF
R1_64 iDFF_9_q_reg:D PNN33_2 4.000000
R2_64 PNN33 PNN33_2 36.935999

C1_297 U167:C 0 0.000127PF
C2_297 n72_4 0 0.000150PF
C3_297 n72_3 0 0.000293PF
C4_297 n72_2 0 0.000293PF
C5_297 U168:Z 0 0.000045PF
R1_297 U168:Z n72_2 4.000000
R2_297 n72_3 n72_2 1.216000
R3_297 n72_3 n72_4 4.000000
R4_297 U167:C n72_4 1.368000

C1_44 PNN105 0 0.002450PF
C2_44 PNN105_6 0 0.002506PF
C3_44 PNN105_5 0 0.000821PF
C4_44 PNN105_4 0 0.000821PF
C5_44 PNN105_3 0 0.000349PF
C6_44 PNN105_2 0 0.000314PF
C7_44 iDFF_27_q_reg:D 0 0.000045PF
R1_44 iDFF_27_q_reg:D PNN105_2 4.000000
R2_44 PNN105_2 PNN105_3 3.800000
R3_44 PNN105_4 PNN105_3 0.152000
R4_44 PNN105_4 PNN105_5 4.864000
R5_44 PNN105_5 PNN105_6 0.152000
R6_44 PNN105_6 PNN105 30.095999

C1_252 clk_r_REG35_S2:Q 0 0.000045PF
C2_252 n31_4 0 0.000128PF
C3_252 n31_3 0 0.000128PF
C4_252 n31_2 0 0.000115PF
C5_252 U292:A 0 0.000093PF
R1_252 n31_2 U292:A 0.760000
R2_252 n31_2 n31_3 4.000000
R3_252 n31_4 n31_3 1.064000
R4_252 n31_4 clk_r_REG35_S2:Q 4.000000

C1_213 U217:Z 0 0.000031PF
C2_213 n150_4 0 0.000053PF
C3_213 n150_3 0 0.000832PF
C4_213 n150_2 0 0.000832PF
C5_213 U216:C 0 0.000045PF
R1_213 U216:C n150_2 4.000000
R2_213 n150_2 n150_3 5.624000
R3_213 n150_3 n150_4 4.000000
R4_213 n150_4 U217:Z 0.304000

C1_126 oDFF_12_q_reg:Q 0 0.000045PF
C2_126 Qout_PNN735_5 0 0.002676PF
C3_126 Qout_PNN735_4 0 0.002676PF
C4_126 Qout_PNN735_3 0 0.000069PF
C5_126 Qout_PNN735_2 0 0.000069PF
C6_126 Qout_PNN735 0 0.000042PF
R1_126 Qout_PNN735 Qout_PNN735_2 4.000000
R2_126 Qout_PNN735_2 Qout_PNN735_3 0.608000
R3_126 Qout_PNN735_3 Qout_PNN735_4 4.000000
R4_126 Qout_PNN735_4 Qout_PNN735_5 32.679999
R5_126 Qout_PNN735_5 oDFF_12_q_reg:Q 4.000000

C1_218 U207:Z 0 0.000045PF
C2_218 n156_5 0 0.000405PF
C3_218 n156_4 0 0.000440PF
C4_218 n156_3 0 0.000575PF
C5_218 n156_2 0 0.000541PF
C6_218 U160:C 0 0.000045PF
R1_218 U160:C n156_2 4.000000
R2_218 n156_2 n156_3 5.776000
R3_218 n156_4 n156_3 0.152000
R4_218 n156_4 n156_5 3.800000
R5_218 n156_5 U207:Z 4.000000

C1_207 U220:C 0 0.000045PF
C2_207 n145_3 0 0.000136PF
C3_207 n145_2 0 0.000136PF
C4_207 U221:Z 0 0.000045PF
R1_207 U221:Z n145_2 4.000000
R2_207 n145_3 n145_2 1.672000
R3_207 n145_3 U220:C 4.000000

C1_124 oDFF_10_q_reg:Q 0 0.000045PF
C2_124 Qout_PNN733_7 0 0.000182PF
C3_124 Qout_PNN733_6 0 0.000217PF
C4_124 Qout_PNN733_5 0 0.002515PF
C5_124 Qout_PNN733_4 0 0.002480PF
C6_124 Qout_PNN733_3 0 0.000104PF
C7_124 Qout_PNN733_2 0 0.000104PF
C8_124 Qout_PNN733 0 0.000042PF
R1_124 Qout_PNN733 Qout_PNN733_2 4.000000
R2_124 Qout_PNN733_3 Qout_PNN733_2 1.064000
R3_124 Qout_PNN733_3 Qout_PNN733_4 4.000000
R4_124 Qout_PNN733_4 Qout_PNN733_5 29.943999
R5_124 Qout_PNN733_6 Qout_PNN733_5 0.152000
R6_124 Qout_PNN733_6 Qout_PNN733_7 2.736000
R7_124 Qout_PNN733_7 oDFF_10_q_reg:Q 4.000000

C1_258 clk_r_REG29_S2:Q 0 0.000031PF
C2_258 n37_4 0 0.000053PF
C3_258 n37_3 0 0.000120PF
C4_258 n37_2 0 0.000120PF
C5_258 U304:A 0 0.000045PF
R1_258 U304:A n37_2 4.000000
R2_258 n37_2 n37_3 1.216000
R3_258 n37_3 n37_4 4.000000
R4_258 clk_r_REG29_S2:Q n37_4 0.304000

C1_209 U226:Z 0 0.000045PF
C2_209 n147_4 0 0.000172PF
C3_209 n147_3 0 0.000172PF
C4_209 n147_2 0 0.000115PF
C5_209 U222:A 0 0.000093PF
R1_209 U222:A n147_2 0.760000
R2_209 n147_2 n147_3 4.000000
R3_209 n147_4 n147_3 1.216000
R4_209 n147_4 U226:Z 4.000000

C1_15 iDFF_37_q_reg:Q 0 0.000045PF
C2_15 INP_PNN133_5 0 0.000112PF
C3_15 INP_PNN133_4 0 0.000147PF
C4_15 INP_PNN133_3 0 0.000189PF
C5_15 INP_PNN133_2 0 0.000155PF
C6_15 U226:A 0 0.000045PF
R1_15 U226:A INP_PNN133_2 4.000000
R2_15 INP_PNN133_3 INP_PNN133_2 0.608000
R3_15 INP_PNN133_4 INP_PNN133_3 0.152000
R4_15 INP_PNN133_5 INP_PNN133_4 0.760000
R5_15 INP_PNN133_5 iDFF_37_q_reg:Q 4.000000

C1_236 U195:Z 0 0.000045PF
C2_236 n172_3 0 0.000105PF
C3_236 n172_2 0 0.000105PF
C4_236 U194:A 0 0.000045PF
R1_236 U194:A n172_2 4.000000
R2_236 n172_3 n172_2 1.064000
R3_236 n172_3 U195:Z 4.000000

C1_228 U213:Z 0 0.000045PF
C2_228 n165_5 0 0.000531PF
C3_228 n165_4 0 0.000565PF
C4_228 n165_3 0 0.000239PF
C5_228 n165_2 0 0.000205PF
C6_228 U212:A 0 0.000045PF
R1_228 U212:A n165_2 4.000000
R2_228 n165_2 n165_3 2.736000
R3_228 n165_4 n165_3 0.152000
R4_228 n165_4 n165_5 4.408000
R5_228 n165_5 U213:Z 4.000000

C1_128 oDFF_14_q_reg:Q 0 0.000045PF
C2_128 Qout_PNN737_5 0 0.002670PF
C3_128 Qout_PNN737_4 0 0.002670PF
C4_128 Qout_PNN737_3 0 0.000069PF
C5_128 Qout_PNN737_2 0 0.000069PF
C6_128 Qout_PNN737 0 0.000042PF
R1_128 Qout_PNN737 Qout_PNN737_2 4.000000
R2_128 Qout_PNN737_2 Qout_PNN737_3 0.608000
R3_128 Qout_PNN737_3 Qout_PNN737_4 4.000000
R4_128 Qout_PNN737_4 Qout_PNN737_5 32.679999
R5_128 Qout_PNN737_5 oDFF_14_q_reg:Q 4.000000

C1_203 U198:Z 0 0.000045PF
C2_203 n140_3 0 0.000107PF
C3_203 n140_2 0 0.000107PF
C4_203 U196:A 0 0.000045PF
R1_203 U196:A n140_2 4.000000
R2_203 n140_3 n140_2 1.520000
R3_203 n140_3 U198:Z 4.000000

C1_229 U255:Z 0 0.000045PF
C2_229 n166_3 0 0.000419PF
C3_229 n166_2 0 0.000419PF
C4_229 U254:A 0 0.000045PF
R1_229 U254:A n166_2 4.000000
R2_229 n166_2 n166_3 5.016000
R3_229 n166_3 U255:Z 4.000000

C1_254 clk_r_REG33_S2:Q 0 0.000045PF
C2_254 n33_4 0 0.000182PF
C3_254 n33_3 0 0.000217PF
C4_254 n33_2 0 0.000086PF
C5_254 U296:A 0 0.000045PF
R1_254 U296:A n33_2 4.000000
R2_254 n33_3 n33_2 0.152000
R3_254 n33_3 n33_4 2.128000
R4_254 n33_4 clk_r_REG33_S2:Q 4.000000

C1_66 PNN41 0 0.000042PF
C2_66 PNN41_5 0 0.000173PF
C3_66 PNN41_4 0 0.000173PF
C4_66 PNN41_3 0 0.002593PF
C5_66 PNN41_2 0 0.002593PF
C6_66 iDFF_11_q_reg:D 0 0.000045PF
R1_66 iDFF_11_q_reg:D PNN41_2 4.000000
R2_66 PNN41_3 PNN41_2 31.311999
R3_66 PNN41_3 PNN41_4 4.000000
R4_66 PNN41_5 PNN41_4 1.976000
R5_66 PNN41_5 PNN41 4.000000

C1_69 PNN5 0 0.002367PF
C2_69 PNN5_6 0 0.002422PF
C3_69 PNN5_5 0 0.001297PF
C4_69 PNN5_4 0 0.001297PF
C5_69 PNN5_3 0 0.000146PF
C6_69 PNN5_2 0 0.000112PF
C7_69 iDFF_2_q_reg:D 0 0.000045PF
R1_69 iDFF_2_q_reg:D PNN5_2 4.000000
R2_69 PNN5_3 PNN5_2 1.368000
R3_69 PNN5_4 PNN5_3 0.152000
R4_69 PNN5_5 PNN5_4 7.904000
R5_69 PNN5_5 PNN5_6 0.152000
R6_69 PNN5 PNN5_6 29.943999

C1_314 U285:Z 0 0.000045PF
C2_314 n88_3 0 0.000160PF
C3_314 n88_2 0 0.000160PF
C4_314 U284:B 0 0.000045PF
R1_314 U284:B n88_2 4.000000
R2_314 n88_3 n88_2 1.824000
R3_314 n88_3 U285:Z 4.000000

C1_102 U284:Z 0 0.000045PF
C2_102 Q_PNN743_4 0 0.000303PF
C3_102 Q_PNN743_3 0 0.000303PF
C4_102 Q_PNN743_2 0 0.000077PF
C5_102 oDFF_20_q_reg:D 0 0.000055PF
R1_102 oDFF_20_q_reg:D Q_PNN743_2 0.608000
R2_102 Q_PNN743_2 Q_PNN743_3 4.000000
R3_102 Q_PNN743_4 Q_PNN743_3 3.648000
R4_102 Q_PNN743_4 U284:Z 4.000000

C1_129 oDFF_15_q_reg:Q 0 0.000045PF
C2_129 Qout_PNN738_5 0 0.003664PF
C3_129 Qout_PNN738_4 0 0.003664PF
C4_129 Qout_PNN738_3 0 0.000046PF
C5_129 Qout_PNN738_2 0 0.000046PF
C6_129 Qout_PNN738 0 0.000042PF
R1_129 Qout_PNN738 Qout_PNN738_2 4.000000
R2_129 Qout_PNN738_3 Qout_PNN738_2 0.304000
R3_129 Qout_PNN738_3 Qout_PNN738_4 4.000000
R4_129 Qout_PNN738_4 Qout_PNN738_5 32.679999
R5_129 Qout_PNN738_5 oDFF_15_q_reg:Q 4.000000

C1_72 PNN61 0 0.000042PF
C2_72 PNN61_9 0 0.000080PF
C3_72 PNN61_8 0 0.000080PF
C4_72 PNN61_7 0 0.000039PF
C5_72 PNN61_6 0 0.000055PF
C6_72 PNN61_5 0 0.000125PF
C7_72 PNN61_4 0 0.000125PF
C8_72 PNN61_3 0 0.002724PF
C9_72 PNN61_2 0 0.002724PF
C10_72 iDFF_16_q_reg:D 0 0.000045PF
R1_72 iDFF_16_q_reg:D PNN61_2 4.000000
R2_72 PNN61_3 PNN61_2 31.159999
R3_72 PNN61_3 PNN61_4 4.000000
R4_72 PNN61_4 PNN61_5 1.368000
R5_72 PNN61_5 PNN61_6 4.000000
R6_72 PNN61_7 PNN61_6 0.152000
R7_72 PNN61_7 PNN61_8 4.000000
R8_72 PNN61_8 PNN61_9 0.760000
R9_72 PNN61_9 PNN61 4.000000

C1_127 oDFF_13_q_reg:Q 0 0.000045PF
C2_127 Qout_PNN736_8 0 0.000121PF
C3_127 Qout_PNN736_7 0 0.000047PF
C4_127 Qout_PNN736_6 0 0.000047PF
C5_127 Qout_PNN736_5 0 0.002776PF
C6_127 Qout_PNN736_4 0 0.002776PF
C7_127 Qout_PNN736_3 0 0.000069PF
C8_127 Qout_PNN736_2 0 0.000069PF
C9_127 Qout_PNN736 0 0.000042PF
R1_127 Qout_PNN736 Qout_PNN736_2 4.000000
R2_127 Qout_PNN736_3 Qout_PNN736_2 0.608000
R3_127 Qout_PNN736_3 Qout_PNN736_4 4.000000
R4_127 Qout_PNN736_4 Qout_PNN736_5 30.703999
R5_127 Qout_PNN736_5 Qout_PNN736_6 4.000000
R6_127 Qout_PNN736_7 Qout_PNN736_6 0.304000
R7_127 Qout_PNN736_7 Qout_PNN736_8 4.000000
R8_127 Qout_PNN736_8 oDFF_13_q_reg:Q 4.000000

C1_70 PNN53 0 0.000042PF
C2_70 PNN53_9 0 0.000115PF
C3_70 PNN53_8 0 0.000115PF
C4_70 PNN53_7 0 0.003389PF
C5_70 PNN53_6 0 0.003389PF
C6_70 PNN53_5 0 0.000062PF
C7_70 PNN53_4 0 0.000062PF
C8_70 PNN53_3 0 0.000374PF
C9_70 PNN53_2 0 0.000374PF
C10_70 iDFF_14_q_reg:D 0 0.000045PF
R1_70 iDFF_14_q_reg:D PNN53_2 4.000000
R2_70 PNN53_3 PNN53_2 2.128000
R3_70 PNN53_3 PNN53_4 4.000000
R4_70 PNN53_5 PNN53_4 0.304000
R5_70 PNN53_5 PNN53_6 4.000000
R6_70 PNN53_7 PNN53_6 30.855999
R7_70 PNN53_7 PNN53_8 4.000000
R8_70 PNN53_8 PNN53_9 1.216000
R9_70 PNN53_9 PNN53 4.000000

C1_266 oDFF_5_q_reg:D 0 0.000045PF
C2_266 n44_7 0 0.000033PF
C3_266 n44_6 0 0.000049PF
C4_266 n44_5 0 0.000056PF
C5_266 n44_4 0 0.000056PF
C6_266 n44_3 0 0.000045PF
C7_266 n44_2 0 0.000045PF
C8_266 clk_r_REG2_S2:Q 0 0.000045PF
R1_266 clk_r_REG2_S2:Q n44_2 4.000000
R2_266 n44_2 n44_3 0.304000
R3_266 n44_3 n44_4 4.000000
R4_266 n44_4 n44_5 0.304000
R5_266 n44_5 n44_6 4.000000
R6_266 n44_6 n44_7 0.152000
R7_266 n44_7 oDFF_5_q_reg:D 4.000000

C1_95 U298:Z 0 0.000045PF
C2_95 Q_PNN736_6 0 0.000121PF
C3_95 Q_PNN736_5 0 0.000143PF
C4_95 Q_PNN736_4 0 0.000143PF
C5_95 Q_PNN736_3 0 0.000069PF
C6_95 Q_PNN736_2 0 0.000069PF
C7_95 oDFF_13_q_reg:D 0 0.000045PF
R1_95 oDFF_13_q_reg:D Q_PNN736_2 4.000000
R2_95 Q_PNN736_3 Q_PNN736_2 0.304000
R3_95 Q_PNN736_3 Q_PNN736_4 4.000000
R4_95 Q_PNN736_4 Q_PNN736_5 1.064000
R5_95 Q_PNN736_5 Q_PNN736_6 4.000000
R6_95 Q_PNN736_6 U298:Z 4.000000

C1_257 U302:A 0 0.000045PF
C2_257 n36_6 0 0.000055PF
C3_257 n36_5 0 0.000071PF
C4_257 n36_4 0 0.000087PF
C5_257 n36_3 0 0.000087PF
C6_257 n36_2 0 0.000121PF
C7_257 clk_r_REG30_S2:Q 0 0.000045PF
R1_257 clk_r_REG30_S2:Q n36_2 4.000000
R2_257 n36_2 n36_3 4.000000
R3_257 n36_3 n36_4 0.608000
R4_257 n36_4 n36_5 4.000000
R5_257 n36_5 n36_6 0.152000
R6_257 n36_6 U302:A 4.000000

C1_93 oDFF_11_q_reg:D 0 0.000045PF
C2_93 Q_PNN734_6 0 0.000033PF
C3_93 Q_PNN734_5 0 0.000049PF
C4_93 Q_PNN734_4 0 0.000057PF
C5_93 Q_PNN734_3 0 0.000057PF
C6_93 Q_PNN734_2 0 0.000121PF
C7_93 U302:Z 0 0.000045PF
R1_93 U302:Z Q_PNN734_2 4.000000
R2_93 Q_PNN734_2 Q_PNN734_3 4.000000
R3_93 Q_PNN734_3 Q_PNN734_4 0.456000
R4_93 Q_PNN734_4 Q_PNN734_5 4.000000
R5_93 Q_PNN734_6 Q_PNN734_5 0.152000
R6_93 Q_PNN734_6 oDFF_11_q_reg:D 4.000000

C1_98 U292:Z 0 0.000045PF
C2_98 Q_PNN739_7 0 0.000142PF
C3_98 Q_PNN739_6 0 0.000142PF
C4_98 Q_PNN739_5 0 0.000183PF
C5_98 Q_PNN739_4 0 0.000183PF
C6_98 Q_PNN739_3 0 0.000043PF
C7_98 Q_PNN739_2 0 0.000043PF
C8_98 oDFF_16_q_reg:D 0 0.000045PF
R1_98 oDFF_16_q_reg:D Q_PNN739_2 4.000000
R2_98 Q_PNN739_2 Q_PNN739_3 0.304000
R3_98 Q_PNN739_3 Q_PNN739_4 4.000000
R4_98 Q_PNN739_4 Q_PNN739_5 1.368000
R5_98 Q_PNN739_5 Q_PNN739_6 4.000000
R6_98 Q_PNN739_6 Q_PNN739_7 1.064000
R7_98 Q_PNN739_7 U292:Z 4.000000

C1_164 U303:Z 0 0.000045PF
C2_164 n100_7 0 0.000083PF
C3_164 n100_6 0 0.000083PF
C4_164 n100_5 0 0.000264PF
C5_164 n100_4 0 0.000264PF
C6_164 n100_3 0 0.000105PF
C7_164 n100_2 0 0.000105PF
C8_164 U302:B 0 0.000045PF
R1_164 U302:B n100_2 4.000000
R2_164 n100_2 n100_3 1.368000
R3_164 n100_3 n100_4 4.000000
R4_164 n100_5 n100_4 3.344000
R5_164 n100_5 n100_6 4.000000
R6_164 n100_6 n100_7 0.456000
R7_164 n100_7 U303:Z 4.000000

C1_87 U315:Z 0 0.000045PF
C2_87 Q_PNN728_6 0 0.000121PF
C3_87 Q_PNN728_5 0 0.000169PF
C4_87 Q_PNN728_4 0 0.000169PF
C5_87 Q_PNN728_3 0 0.000129PF
C6_87 Q_PNN728_2 0 0.000129PF
C7_87 clk_r_REG2_S2:D 0 0.000045PF
R1_87 clk_r_REG2_S2:D Q_PNN728_2 4.000000
R2_87 Q_PNN728_2 Q_PNN728_3 1.368000
R3_87 Q_PNN728_3 Q_PNN728_4 4.000000
R4_87 Q_PNN728_4 Q_PNN728_5 1.824000
R5_87 Q_PNN728_5 Q_PNN728_6 4.000000
R6_87 Q_PNN728_6 U315:Z 4.000000

C1_96 oDFF_14_q_reg:D 0 0.000045PF
C2_96 Q_PNN737_5 0 0.000121PF
C3_96 Q_PNN737_4 0 0.000058PF
C4_96 Q_PNN737_3 0 0.000058PF
C5_96 Q_PNN737_2 0 0.000121PF
C6_96 U296:Z 0 0.000045PF
R1_96 U296:Z Q_PNN737_2 4.000000
R2_96 Q_PNN737_2 Q_PNN737_3 4.000000
R3_96 Q_PNN737_4 Q_PNN737_3 0.456000
R4_96 Q_PNN737_4 Q_PNN737_5 4.000000
R5_96 Q_PNN737_5 oDFF_14_q_reg:D 4.000000

C1_320 U292:B 0 0.000045PF
C2_320 n93_5 0 0.000121PF
C3_320 n93_4 0 0.000125PF
C4_320 n93_3 0 0.000125PF
C5_320 n93_2 0 0.000121PF
C6_320 U293:Z 0 0.000045PF
R1_320 U293:Z n93_2 4.000000
R2_320 n93_2 n93_3 4.000000
R3_320 n93_4 n93_3 1.064000
R4_320 n93_4 n93_5 4.000000
R5_320 n93_5 U292:B 4.000000

C1_323 U297:Z 0 0.000045PF
C2_323 n96_6 0 0.000218PF
C3_323 n96_5 0 0.000218PF
C4_323 n96_4 0 0.000045PF
C5_323 n96_3 0 0.000045PF
C6_323 n96_2 0 0.000121PF
C7_323 U296:B 0 0.000045PF
R1_323 U296:B n96_2 4.000000
R2_323 n96_2 n96_3 4.000000
R3_323 n96_3 n96_4 0.304000
R4_323 n96_4 n96_5 4.000000
R5_323 n96_5 n96_6 1.824000
R6_323 n96_6 U297:Z 4.000000

C1_171 U316:Z 0 0.000045PF
C2_171 n107_7 0 0.000162PF
C3_171 n107_6 0 0.000162PF
C4_171 n107_5 0 0.000174PF
C5_171 n107_4 0 0.000174PF
C6_171 n107_3 0 0.000045PF
C7_171 n107_2 0 0.000045PF
C8_171 U315:B 0 0.000045PF
R1_171 U315:B n107_2 4.000000
R2_171 n107_2 n107_3 0.304000
R3_171 n107_3 n107_4 4.000000
R4_171 n107_4 n107_5 1.064000
R5_171 n107_5 n107_6 4.000000
R6_171 n107_6 n107_7 1.672000
R7_171 n107_7 U316:Z 4.000000

C1_160 iDFF_5_q_reg:QN 0 0.000045PF
C2_160 c0_n9_12 0 0.000121PF
C3_160 c0_n9_10 0 0.000341PF
C4_160 c0_n9_8 0 0.000112PF
C5_160 c0_n9_6 0 0.000244PF
C6_160 c0_n9_4 0 0.000244PF
C7_160 U315:A 0 0.000045PF
C8_160 c0_n9_15 0 0.000034PF
C9_160 c0_n9_13 0 0.000050PF
C10_160 c0_n9_11 0 0.000248PF
C11_160 U251:A 0 0.000045PF
C12_160 c0_n9_7 0 0.000151PF
C13_160 c0_n9_5 0 0.000186PF
C14_160 c0_n9_3 0 0.000234PF
C15_160 c0_n9_2 0 0.000200PF
C16_160 U239:A 0 0.000090PF
R1_160 U239:A c0_n9_2 4.000000
R2_160 c0_n9_2 c0_n9_3 1.064000
R3_160 U239:A c0_n9_4 4.000000
R4_160 c0_n9_5 c0_n9_3 0.152000
R5_160 c0_n9_6 c0_n9_4 3.192000
R6_160 c0_n9_5 c0_n9_7 1.064000
R7_160 c0_n9_6 c0_n9_8 4.000000
R8_160 c0_n9_7 U251:A 4.000000
R9_160 c0_n9_10 c0_n9_8 2.128000
R10_160 c0_n9_11 c0_n9_10 3.192000
R11_160 c0_n9_10 c0_n9_12 4.000000
R12_160 c0_n9_11 c0_n9_13 4.000000
R13_160 c0_n9_12 iDFF_5_q_reg:QN 4.000000
R14_160 c0_n9_13 c0_n9_15 0.152000
R15_160 c0_n9_15 U315:A 4.000000

C1_94 U300:Z 0 0.000045PF
C2_94 Q_PNN735_7 0 0.000036PF
C3_94 Q_PNN735_6 0 0.000052PF
C4_94 Q_PNN735_5 0 0.000382PF
C5_94 Q_PNN735_4 0 0.000382PF
C6_94 Q_PNN735_3 0 0.000393PF
C7_94 Q_PNN735_2 0 0.000393PF
C8_94 oDFF_12_q_reg:D 0 0.000045PF
R1_94 oDFF_12_q_reg:D Q_PNN735_2 4.000000
R2_94 Q_PNN735_2 Q_PNN735_3 1.672000
R3_94 Q_PNN735_3 Q_PNN735_4 4.000000
R4_94 Q_PNN735_4 Q_PNN735_5 1.824000
R5_94 Q_PNN735_5 Q_PNN735_6 4.000000
R6_94 Q_PNN735_6 Q_PNN735_7 0.152000
R7_94 Q_PNN735_7 U300:Z 4.000000

C1_92 U304:Z 0 0.000045PF
C2_92 Q_PNN733_7 0 0.000032PF
C3_92 Q_PNN733_6 0 0.000049PF
C4_92 Q_PNN733_5 0 0.000114PF
C5_92 Q_PNN733_4 0 0.000114PF
C6_92 Q_PNN733_3 0 0.000153PF
C7_92 Q_PNN733_2 0 0.000153PF
C8_92 oDFF_10_q_reg:D 0 0.000045PF
R1_92 oDFF_10_q_reg:D Q_PNN733_2 4.000000
R2_92 Q_PNN733_2 Q_PNN733_3 1.672000
R3_92 Q_PNN733_3 Q_PNN733_4 4.000000
R4_92 Q_PNN733_5 Q_PNN733_4 0.912000
R5_92 Q_PNN733_5 Q_PNN733_6 4.000000
R6_92 Q_PNN733_6 Q_PNN733_7 0.152000
R7_92 Q_PNN733_7 U304:Z 4.000000

C1_97 U294:Z 0 0.000045PF
C2_97 Q_PNN738_7 0 0.000032PF
C3_97 Q_PNN738_6 0 0.000049PF
C4_97 Q_PNN738_5 0 0.000063PF
C5_97 Q_PNN738_4 0 0.000063PF
C6_97 Q_PNN738_3 0 0.000148PF
C7_97 Q_PNN738_2 0 0.000148PF
C8_97 oDFF_15_q_reg:D 0 0.000045PF
R1_97 oDFF_15_q_reg:D Q_PNN738_2 4.000000
R2_97 Q_PNN738_2 Q_PNN738_3 1.672000
R3_97 Q_PNN738_3 Q_PNN738_4 4.000000
R4_97 Q_PNN738_5 Q_PNN738_4 0.760000
R5_97 Q_PNN738_5 Q_PNN738_6 4.000000
R6_97 Q_PNN738_6 Q_PNN738_7 0.152000
R7_97 Q_PNN738_7 U294:Z 4.000000

C1_325 U301:Z 0 0.000045PF
C2_325 n98_7 0 0.000039PF
C3_325 n98_6 0 0.000055PF
C4_325 n98_5 0 0.000454PF
C5_325 n98_4 0 0.000454PF
C6_325 n98_3 0 0.000050PF
C7_325 n98_2 0 0.000034PF
C8_325 U300:B 0 0.000045PF
R1_325 U300:B n98_2 4.000000
R2_325 n98_3 n98_2 0.152000
R3_325 n98_3 n98_4 4.000000
R4_325 n98_5 n98_4 3.496000
R5_325 n98_5 n98_6 4.000000
R6_325 n98_6 n98_7 0.152000
R7_325 n98_7 U301:Z 4.000000

C1_166 U307:Z 0 0.000045PF
C2_166 n102_6 0 0.000121PF
C3_166 n102_5 0 0.000049PF
C4_166 n102_4 0 0.000049PF
C5_166 n102_3 0 0.000164PF
C6_166 n102_2 0 0.000164PF
C7_166 U306:B 0 0.000045PF
R1_166 U306:B n102_2 4.000000
R2_166 n102_3 n102_2 2.128000
R3_166 n102_3 n102_4 4.000000
R4_166 n102_4 n102_5 0.456000
R5_166 n102_5 n102_6 4.000000
R6_166 n102_6 U307:Z 4.000000

C1_165 U304:B 0 0.000045PF
C2_165 n101_5 0 0.000121PF
C3_165 n101_4 0 0.000083PF
C4_165 n101_3 0 0.000083PF
C5_165 n101_2 0 0.000121PF
C6_165 U305:Z 0 0.000045PF
R1_165 U305:Z n101_2 4.000000
R2_165 n101_2 n101_3 4.000000
R3_165 n101_4 n101_3 0.608000
R4_165 n101_4 n101_5 4.000000
R5_165 n101_5 U304:B 4.000000

C1_322 U295:Z 0 0.000045PF
C2_322 n95_5 0 0.000121PF
C3_322 n95_4 0 0.000664PF
C4_322 n95_3 0 0.000664PF
C5_322 n95_2 0 0.000121PF
C6_322 U294:B 0 0.000045PF
R1_322 U294:B n95_2 4.000000
R2_322 n95_2 n95_3 4.000000
R3_322 n95_4 n95_3 6.688000
R4_322 n95_4 n95_5 4.000000
R5_322 n95_5 U295:Z 4.000000

C1_90 U234:Z 0 0.000045PF
C2_90 Q_PNN731_5 0 0.000121PF
C3_90 Q_PNN731_4 0 0.000236PF
C4_90 Q_PNN731_3 0 0.000236PF
C5_90 Q_PNN731_2 0 0.000121PF
C6_90 clk_r_REG7_S2:D 0 0.000045PF
R1_90 clk_r_REG7_S2:D Q_PNN731_2 4.000000
R2_90 Q_PNN731_2 Q_PNN731_3 4.000000
R3_90 Q_PNN731_3 Q_PNN731_4 2.736000
R4_90 Q_PNN731_4 Q_PNN731_5 4.000000
R5_90 Q_PNN731_5 U234:Z 4.000000

C1_202 clk_r_REG0_S2:Q 0 0.000045PF
C2_202 n14_8 0 0.000121PF
C3_202 n14_7 0 0.000089PF
C4_202 n14_6 0 0.000089PF
C5_202 n14_5 0 0.000121PF
C6_202 U307:A 0 0.000090PF
C7_202 n14_3 0 0.000268PF
C8_202 n14_2 0 0.000268PF
C9_202 U299:A 0 0.000045PF
R1_202 U299:A n14_2 4.000000
R2_202 n14_2 n14_3 2.128000
R3_202 n14_3 U307:A 4.000000
R4_202 U307:A n14_5 4.000000
R5_202 n14_5 n14_6 4.000000
R6_202 n14_7 n14_6 1.064000
R7_202 n14_7 n14_8 4.000000
R8_202 n14_8 clk_r_REG0_S2:Q 4.000000

C1_283 U293:A 0 0.000045PF
C2_283 n6_10 0 0.000122PF
C3_283 n6_8 0 0.000157PF
C4_283 n6_6 0 0.000105PF
C5_283 n6_4 0 0.000070PF
C6_283 clk_r_REG23_S2:Q 0 0.000045PF
C7_283 n6_7 0 0.000121PF
C8_283 n6_5 0 0.001073PF
C9_283 n6_3 0 0.001073PF
C10_283 n6_2 0 0.000121PF
C11_283 U301:A 0 0.000090PF
R1_283 U301:A n6_2 4.000000
R2_283 n6_2 n6_3 4.000000
R3_283 U301:A n6_4 4.000000
R4_283 n6_5 n6_3 4.712000
R5_283 n6_6 n6_4 0.912000
R6_283 n6_5 n6_7 4.000000
R7_283 n6_8 n6_6 0.152000
R8_283 n6_7 clk_r_REG23_S2:Q 4.000000
R9_283 n6_10 n6_8 1.216000
R10_283 n6_10 U293:A 4.000000

C1_272 clk_r_REG19_S2:Q 0 0.000045PF
C2_272 n5_8 0 0.000125PF
C3_272 n5_5 0 0.000125PF
C4_272 n5_2 0 0.000519PF
C5_272 n5_4 0 0.000242PF
C6_272 n5_7 0 0.000121PF
C7_272 U297:A 0 0.000045PF
C8_272 U305:A 0 0.000045PF
C9_272 n5_3 0 0.000121PF
C10_272 n5_1 0 0.000295PF
R1_272 n5_1 n5_2 1.216000
R2_272 n5_1 n5_3 4.000000
R3_272 n5_2 n5_4 1.672000
R4_272 n5_2 n5_5 4.000000
R5_272 n5_3 U305:A 4.000000
R6_272 n5_4 n5_7 4.000000
R7_272 n5_5 n5_8 1.216000
R8_272 n5_7 U297:A 4.000000
R9_272 n5_8 clk_r_REG19_S2:Q 4.000000

C1_253 clk_r_REG34_S2:Q 0 0.000045PF
C2_253 n32_6 0 0.000121PF
C3_253 n32_5 0 0.000340PF
C4_253 n32_4 0 0.000340PF
C5_253 n32_3 0 0.000049PF
C6_253 n32_2 0 0.000032PF
C7_253 U294:A 0 0.000045PF
R1_253 U294:A n32_2 4.000000
R2_253 n32_3 n32_2 0.152000
R3_253 n32_3 n32_4 4.000000
R4_253 n32_5 n32_4 3.344000
R5_253 n32_5 n32_6 4.000000
R6_253 n32_6 clk_r_REG34_S2:Q 4.000000

C1_256 U300:A 0 0.000045PF
C2_256 n35_6 0 0.000121PF
C3_256 n35_5 0 0.000298PF
C4_256 n35_4 0 0.000298PF
C5_256 n35_3 0 0.000050PF
C6_256 n35_2 0 0.000033PF
C7_256 clk_r_REG31_S2:Q 0 0.000045PF
R1_256 clk_r_REG31_S2:Q n35_2 4.000000
R2_256 n35_2 n35_3 0.152000
R3_256 n35_3 n35_4 4.000000
R4_256 n35_4 n35_5 0.760000
R5_256 n35_5 n35_6 4.000000
R6_256 n35_6 U300:A 4.000000

C1_294 clk_r_REG20_S2:Q 0 0.000045PF
C2_294 n7_10 0 0.000255PF
C3_294 n7_9 0 0.000255PF
C4_294 n7_8 0 0.000182PF
C5_294 n7_7 0 0.000182PF
C6_294 n7_6 0 0.000052PF
C7_294 n7_5 0 0.000035PF
C8_294 U295:A 0 0.000090PF
C9_294 n7_3 0 0.000293PF
C10_294 n7_2 0 0.000293PF
C11_294 U303:A 0 0.000045PF
R1_294 U303:A n7_2 4.000000
R2_294 n7_2 n7_3 2.128000
R3_294 n7_3 U295:A 4.000000
R4_294 U295:A n7_5 4.000000
R5_294 n7_5 n7_6 0.152000
R6_294 n7_6 n7_7 4.000000
R7_294 n7_7 n7_8 1.368000
R8_294 n7_8 n7_9 4.000000
R9_294 n7_9 n7_10 1.064000
R10_294 n7_10 clk_r_REG20_S2:Q 4.000000

C1_223 U253:Z 0 0.000045PF
C2_223 n160_6 0 0.000222PF
C3_223 n160_5 0 0.000222PF
C4_223 n160_4 0 0.000178PF
C5_223 n160_3 0 0.000178PF
C6_223 n160_2 0 0.000121PF
C7_223 U252:A 0 0.000095PF
R1_223 U252:A n160_2 2.000000
R2_223 n160_2 n160_3 4.000000
R3_223 n160_3 n160_4 1.976000
R4_223 n160_4 n160_5 4.000000
R5_223 n160_6 n160_5 1.064000
R6_223 n160_6 U253:Z 4.000000

C1_269 clk_r_REG9_S2:Q 0 0.000045PF
C2_269 n47_7 0 0.000034PF
C3_269 n47_6 0 0.000050PF
C4_269 n47_5 0 0.000110PF
C5_269 n47_4 0 0.000110PF
C6_269 n47_3 0 0.000040PF
C7_269 n47_2 0 0.000040PF
C8_269 oDFF_2_q_reg:D 0 0.000045PF
R1_269 oDFF_2_q_reg:D n47_2 4.000000
R2_269 n47_3 n47_2 0.304000
R3_269 n47_3 n47_4 4.000000
R4_269 n47_5 n47_4 0.760000
R5_269 n47_5 n47_6 4.000000
R6_269 n47_6 n47_7 0.152000
R7_269 n47_7 clk_r_REG9_S2:Q 4.000000

C1_259 U306:A 0 0.000045PF
C2_259 n38_6 0 0.000076PF
C3_259 n38_5 0 0.000093PF
C4_259 n38_4 0 0.000182PF
C5_259 n38_3 0 0.000182PF
C6_259 n38_2 0 0.000121PF
C7_259 clk_r_REG26_S2:Q 0 0.000045PF
R1_259 clk_r_REG26_S2:Q n38_2 4.000000
R2_259 n38_2 n38_3 4.000000
R3_259 n38_4 n38_3 2.128000
R4_259 n38_4 n38_5 4.000000
R5_259 n38_6 n38_5 0.152000
R6_259 n38_6 U306:A 4.000000

C1_91 oDFF_9_q_reg:D 0 0.000045PF
C2_91 Q_PNN732_5 0 0.000121PF
C3_91 Q_PNN732_4 0 0.000095PF
C4_91 Q_PNN732_3 0 0.000095PF
C5_91 Q_PNN732_2 0 0.000121PF
C6_91 U306:Z 0 0.000045PF
R1_91 U306:Z Q_PNN732_2 4.000000
R2_91 Q_PNN732_2 Q_PNN732_3 4.000000
R3_91 Q_PNN732_4 Q_PNN732_3 0.912000
R4_91 Q_PNN732_4 Q_PNN732_5 4.000000
R5_91 Q_PNN732_5 oDFF_9_q_reg:D 4.000000

C1_116 oDFF_2_q_reg:Q 0 0.000045PF
C2_116 Qout_PNN725_7 0 0.000044PF
C3_116 Qout_PNN725_6 0 0.000044PF
C4_116 Qout_PNN725_5 0 0.002436PF
C5_116 Qout_PNN725_4 0 0.002436PF
C6_116 Qout_PNN725_3 0 0.000044PF
C7_116 Qout_PNN725_2 0 0.000044PF
C8_116 Qout_PNN725 0 0.000042PF
R1_116 Qout_PNN725 Qout_PNN725_2 4.000000
R2_116 Qout_PNN725_2 Qout_PNN725_3 0.304000
R3_116 Qout_PNN725_3 Qout_PNN725_4 4.000000
R4_116 Qout_PNN725_5 Qout_PNN725_4 30.551999
R5_116 Qout_PNN725_5 Qout_PNN725_6 4.000000
R6_116 Qout_PNN725_7 Qout_PNN725_6 0.304000
R7_116 Qout_PNN725_7 oDFF_2_q_reg:Q 4.000000

C1_27 U252:C 0 0.000045PF
C2_27 INP_PNN49_11 0 0.000034PF
C3_27 INP_PNN49_9 0 0.000096PF
C4_27 INP_PNN49_7 0 0.001241PF
C5_27 INP_PNN49_4 0 0.001241PF
C6_27 INP_PNN49_2 0 0.000447PF
C7_27 U239:B 0 0.000045PF
C8_27 clk_r_REG32_S2:D 0 0.000045PF
C9_27 INP_PNN49_19 0 0.000046PF
C10_27 INP_PNN49_18 0 0.000046PF
C11_27 INP_PNN49_17 0 0.000075PF
C12_27 INP_PNN49_16 0 0.000075PF
C13_27 INP_PNN49_15 0 0.000106PF
C14_27 INP_PNN49_14 0 0.000106PF
C15_27 iDFF_13_q_reg:Q 0 0.000090PF
C16_27 INP_PNN49_10 0 0.000145PF
C17_27 INP_PNN49_8 0 0.000145PF
C18_27 INP_PNN49_6 0 0.000206PF
C19_27 INP_PNN49_3 0 0.000206PF
C20_27 INP_PNN49_1 0 0.000447PF
R1_27 INP_PNN49_1 INP_PNN49_2 2.128000
R2_27 INP_PNN49_1 INP_PNN49_3 4.000000
R3_27 INP_PNN49_2 INP_PNN49_4 4.000000
R4_27 INP_PNN49_2 U239:B 4.000000
R5_27 INP_PNN49_3 INP_PNN49_6 2.128000
R6_27 INP_PNN49_4 INP_PNN49_7 9.880000
R7_27 INP_PNN49_6 INP_PNN49_8 4.000000
R8_27 INP_PNN49_7 INP_PNN49_9 4.000000
R9_27 INP_PNN49_10 INP_PNN49_8 1.520000
R10_27 INP_PNN49_11 INP_PNN49_9 0.152000
R11_27 INP_PNN49_10 iDFF_13_q_reg:Q 4.000000
R12_27 INP_PNN49_11 U252:C 4.000000
R13_27 iDFF_13_q_reg:Q INP_PNN49_14 4.000000
R14_27 INP_PNN49_15 INP_PNN49_14 1.064000
R15_27 INP_PNN49_15 INP_PNN49_16 4.000000
R16_27 INP_PNN49_17 INP_PNN49_16 0.456000
R17_27 INP_PNN49_17 INP_PNN49_18 4.000000
R18_27 INP_PNN49_19 INP_PNN49_18 0.304000
R19_27 INP_PNN49_19 clk_r_REG32_S2:D 4.000000

C1_177 U233:Z 0 0.000045PF
C2_177 n112_6 0 0.000229PF
C3_177 n112_5 0 0.000229PF
C4_177 n112_4 0 0.000288PF
C5_177 n112_3 0 0.000288PF
C6_177 n112_2 0 0.000121PF
C7_177 U232:B 0 0.000045PF
R1_177 U232:B n112_2 4.000000
R2_177 n112_2 n112_3 4.000000
R3_177 n112_4 n112_3 2.736000
R4_177 n112_4 n112_5 4.000000
R5_177 n112_5 n112_6 1.824000
R6_177 n112_6 U233:Z 4.000000

C1_84 clk_r_REG9_S2:D 0 0.000045PF
C2_84 Q_PNN725_6 0 0.000034PF
C3_84 Q_PNN725_5 0 0.000050PF
C4_84 Q_PNN725_4 0 0.000128PF
C5_84 Q_PNN725_3 0 0.000128PF
C6_84 Q_PNN725_2 0 0.000121PF
C7_84 U232:Z 0 0.000045PF
R1_84 U232:Z Q_PNN725_2 4.000000
R2_84 Q_PNN725_2 Q_PNN725_3 4.000000
R3_84 Q_PNN725_3 Q_PNN725_4 0.912000
R4_84 Q_PNN725_4 Q_PNN725_5 4.000000
R5_84 Q_PNN725_6 Q_PNN725_5 0.152000
R6_84 Q_PNN725_6 clk_r_REG9_S2:D 4.000000

C1_274 clk_r_REG1_S2:Q 0 0.000045PF
C2_274 n51_7 0 0.000123PF
C3_274 n51_6 0 0.000123PF
C4_274 n51_5 0 0.000075PF
C5_274 n51_4 0 0.000075PF
C6_274 n51_3 0 0.000047PF
C7_274 n51_2 0 0.000047PF
C8_274 oDFF_1_q_reg:D 0 0.000045PF
R1_274 oDFF_1_q_reg:D n51_2 4.000000
R2_274 n51_2 n51_3 0.456000
R3_274 n51_3 n51_4 4.000000
R4_274 n51_4 n51_5 0.456000
R5_274 n51_5 n51_6 4.000000
R6_274 n51_6 n51_7 1.368000
R7_274 n51_7 clk_r_REG1_S2:Q 4.000000

C1_29 iDFF_14_q_reg:Q 0 0.000045PF
C2_29 INP_PNN53_12 0 0.000424PF
C3_29 INP_PNN53_8 0 0.000424PF
C4_29 INP_PNN53_4 0 0.000354PF
C5_29 INP_PNN53_7 0 0.000187PF
C6_29 INP_PNN53_11 0 0.000121PF
C7_29 U252:B 0 0.000045PF
C8_29 U195:A 0 0.000045PF
C9_29 INP_PNN53_9 0 0.000110PF
C10_29 INP_PNN53_5 0 0.000110PF
C11_29 INP_PNN53_2 0 0.000306PF
C12_29 clk_r_REG33_S2:D 0 0.000045PF
C13_29 INP_PNN53_6 0 0.000169PF
C14_29 INP_PNN53_3 0 0.000169PF
C15_29 INP_PNN53_1 0 0.000139PF
R1_29 INP_PNN53_2 INP_PNN53_1 1.368000
R2_29 INP_PNN53_1 INP_PNN53_3 4.000000
R3_29 INP_PNN53_4 INP_PNN53_2 1.976000
R4_29 INP_PNN53_2 INP_PNN53_5 4.000000
R5_29 INP_PNN53_6 INP_PNN53_3 2.280000
R6_29 INP_PNN53_7 INP_PNN53_4 1.976000
R7_29 INP_PNN53_4 INP_PNN53_8 4.000000
R8_29 INP_PNN53_5 INP_PNN53_9 1.064000
R9_29 INP_PNN53_6 clk_r_REG33_S2:D 4.000000
R10_29 INP_PNN53_7 INP_PNN53_11 4.000000
R11_29 INP_PNN53_12 INP_PNN53_8 4.104000
R12_29 INP_PNN53_9 U195:A 4.000000
R13_29 INP_PNN53_11 U252:B 4.000000
R14_29 INP_PNN53_12 iDFF_14_q_reg:Q 4.000000

C1_22 U251:B 0 0.000045PF
C2_22 INP_PNN29_8 0 0.000057PF
C3_22 INP_PNN29_5 0 0.000057PF
C4_22 INP_PNN29_2 0 0.001428PF
C5_22 INP_PNN29_4 0 0.000926PF
C6_22 INP_PNN29_7 0 0.000050PF
C7_22 INP_PNN29_10 0 0.000034PF
C8_22 U192:B 0 0.000045PF
C9_22 U234:A 0 0.000056PF
C10_22 INP_PNN29_15 0 0.000078PF
C11_22 INP_PNN29_14 0 0.000100PF
C12_22 INP_PNN29_13 0 0.000100PF
C13_22 iDFF_8_q_reg:Q 0 0.000090PF
C14_22 INP_PNN29_6 0 0.000121PF
C15_22 INP_PNN29_3 0 0.000121PF
C16_22 INP_PNN29_1 0 0.000520PF
R1_22 INP_PNN29_1 INP_PNN29_2 5.776000
R2_22 INP_PNN29_1 INP_PNN29_3 4.000000
R3_22 INP_PNN29_2 INP_PNN29_4 5.472000
R4_22 INP_PNN29_2 INP_PNN29_5 4.000000
R5_22 INP_PNN29_6 INP_PNN29_3 1.216000
R6_22 INP_PNN29_4 INP_PNN29_7 4.000000
R7_22 INP_PNN29_5 INP_PNN29_8 0.304000
R8_22 INP_PNN29_6 iDFF_8_q_reg:Q 4.000000
R9_22 INP_PNN29_10 INP_PNN29_7 0.152000
R10_22 INP_PNN29_8 U251:B 4.000000
R11_22 INP_PNN29_10 U192:B 4.000000
R12_22 iDFF_8_q_reg:Q INP_PNN29_13 4.000000
R13_22 INP_PNN29_14 INP_PNN29_13 1.064000
R14_22 INP_PNN29_14 INP_PNN29_15 4.000000
R15_22 INP_PNN29_15 U234:A 0.456000

C1_117 oDFF_3_q_reg:Q 0 0.000045PF
C2_117 Qout_PNN726_7 0 0.000044PF
C3_117 Qout_PNN726_6 0 0.000044PF
C4_117 Qout_PNN726_5 0 0.003194PF
C5_117 Qout_PNN726_4 0 0.003194PF
C6_117 Qout_PNN726_3 0 0.000067PF
C7_117 Qout_PNN726_2 0 0.000067PF
C8_117 Qout_PNN726 0 0.000042PF
R1_117 Qout_PNN726 Qout_PNN726_2 4.000000
R2_117 Qout_PNN726_3 Qout_PNN726_2 0.608000
R3_117 Qout_PNN726_3 Qout_PNN726_4 4.000000
R4_117 Qout_PNN726_5 Qout_PNN726_4 30.551999
R5_117 Qout_PNN726_5 Qout_PNN726_6 4.000000
R6_117 Qout_PNN726_7 Qout_PNN726_6 0.304000
R7_117 Qout_PNN726_7 oDFF_3_q_reg:Q 4.000000

C1_26 clk_r_REG31_S2:D 0 0.000045PF
C2_26 INP_PNN45_17 0 0.000073PF
C3_26 INP_PNN45_16 0 0.000073PF
C4_26 INP_PNN45_15 0 0.000077PF
C5_26 INP_PNN45_14 0 0.000077PF
C6_26 INP_PNN45_13 0 0.000049PF
C7_26 INP_PNN45_12 0 0.000033PF
C8_26 iDFF_12_q_reg:Q 0 0.000090PF
C9_26 INP_PNN45_8 0 0.000172PF
C10_26 INP_PNN45_5 0 0.000172PF
C11_26 INP_PNN45_2 0 0.000149PF
C12_26 INP_PNN45_4 0 0.000078PF
C13_26 INP_PNN45_7 0 0.000121PF
C14_26 U193:B 0 0.000045PF
C15_26 U191:A 0 0.000045PF
C16_26 INP_PNN45_6 0 0.000119PF
C17_26 INP_PNN45_3 0 0.000119PF
C18_26 INP_PNN45_1 0 0.000090PF
R1_26 INP_PNN45_2 INP_PNN45_1 0.760000
R2_26 INP_PNN45_1 INP_PNN45_3 4.000000
R3_26 INP_PNN45_4 INP_PNN45_2 0.912000
R4_26 INP_PNN45_2 INP_PNN45_5 4.000000
R5_26 INP_PNN45_3 INP_PNN45_6 1.824000
R6_26 INP_PNN45_4 INP_PNN45_7 4.000000
R7_26 INP_PNN45_8 INP_PNN45_5 1.672000
R8_26 INP_PNN45_6 U191:A 4.000000
R9_26 INP_PNN45_7 U193:B 4.000000
R10_26 INP_PNN45_8 iDFF_12_q_reg:Q 4.000000
R11_26 iDFF_12_q_reg:Q INP_PNN45_12 4.000000
R12_26 INP_PNN45_13 INP_PNN45_12 0.152000
R13_26 INP_PNN45_13 INP_PNN45_14 4.000000
R14_26 INP_PNN45_14 INP_PNN45_15 0.456000
R15_26 INP_PNN45_15 INP_PNN45_16 4.000000
R16_26 INP_PNN45_17 INP_PNN45_16 1.216000
R17_26 INP_PNN45_17 clk_r_REG31_S2:D 4.000000

C1_28 U232:A 0 0.000045PF
C2_28 INP_PNN5_15 0 0.000057PF
C3_28 INP_PNN5_14 0 0.000091PF
C4_28 INP_PNN5_13 0 0.000127PF
C5_28 INP_PNN5_12 0 0.000093PF
C6_28 iDFF_2_q_reg:Q 0 0.000090PF
C7_28 INP_PNN5_9 0 0.000033PF
C8_28 INP_PNN5_7 0 0.000049PF
C9_28 INP_PNN5_4 0 0.000956PF
C10_28 INP_PNN5_2 0 0.001339PF
C11_28 INP_PNN5_5 0 0.000152PF
C12_28 INP_PNN5_8 0 0.000152PF
C13_28 U249:B 0 0.000045PF
C14_28 U195:B 0 0.000045PF
C15_28 INP_PNN5_3 0 0.000121PF
C16_28 INP_PNN5_1 0 0.000402PF
R1_28 INP_PNN5_1 INP_PNN5_2 1.672000
R2_28 INP_PNN5_1 INP_PNN5_3 4.000000
R3_28 INP_PNN5_2 INP_PNN5_4 6.536000
R4_28 INP_PNN5_2 INP_PNN5_5 4.000000
R5_28 INP_PNN5_3 U195:B 4.000000
R6_28 INP_PNN5_4 INP_PNN5_7 4.000000
R7_28 INP_PNN5_5 INP_PNN5_8 1.824000
R8_28 INP_PNN5_7 INP_PNN5_9 0.152000
R9_28 INP_PNN5_8 U249:B 4.000000
R10_28 INP_PNN5_9 iDFF_2_q_reg:Q 4.000000
R11_28 iDFF_2_q_reg:Q INP_PNN5_12 4.000000
R12_28 INP_PNN5_13 INP_PNN5_12 0.912000
R13_28 INP_PNN5_13 INP_PNN5_14 0.152000
R14_28 INP_PNN5_15 INP_PNN5_14 0.760000
R15_28 INP_PNN5_15 U232:A 4.000000

C1_83 U246:Z 0 0.000045PF
C2_83 Q_PNN724_6 0 0.000121PF
C3_83 Q_PNN724_5 0 0.000687PF
C4_83 Q_PNN724_4 0 0.000687PF
C5_83 Q_PNN724_3 0 0.000050PF
C6_83 Q_PNN724_2 0 0.000034PF
C7_83 clk_r_REG1_S2:D 0 0.000045PF
R1_83 clk_r_REG1_S2:D Q_PNN724_2 4.000000
R2_83 Q_PNN724_2 Q_PNN724_3 0.152000
R3_83 Q_PNN724_3 Q_PNN724_4 4.000000
R4_83 Q_PNN724_4 Q_PNN724_5 4.408000
R5_83 Q_PNN724_5 Q_PNN724_6 4.000000
R6_83 Q_PNN724_6 U246:Z 4.000000

C1_235 U193:Z 0 0.000045PF
C2_235 n171_5 0 0.000121PF
C3_235 n171_4 0 0.000119PF
C4_235 n171_3 0 0.000119PF
C5_235 n171_2 0 0.000121PF
C6_235 U192:A 0 0.000045PF
R1_235 U192:A n171_2 4.000000
R2_235 n171_2 n171_3 4.000000
R3_235 n171_3 n171_4 1.824000
R4_235 n171_4 n171_5 4.000000
R5_235 n171_5 U193:Z 4.000000

C1_80 PNN9 0 0.001072PF
C2_80 PNN9_6 0 0.001128PF
C3_80 PNN9_5 0 0.002346PF
C4_80 PNN9_4 0 0.002312PF
C5_80 PNN9_3 0 0.000050PF
C6_80 PNN9_2 0 0.000034PF
C7_80 iDFF_3_q_reg:D 0 0.000045PF
R1_80 iDFF_3_q_reg:D PNN9_2 4.000000
R2_80 PNN9_2 PNN9_3 0.152000
R3_80 PNN9_3 PNN9_4 4.000000
R4_80 PNN9_4 PNN9_5 24.167999
R5_80 PNN9_6 PNN9_5 0.152000
R6_80 PNN9_6 PNN9 9.120000

C1_2 U248:C 0 0.000045PF
C2_2 INP_PNN1_9 0 0.000233PF
C3_2 INP_PNN1_7 0 0.000233PF
C4_2 INP_PNN1_4 0 0.000094PF
C5_2 INP_PNN1_2 0 0.000593PF
C6_2 INP_PNN1_5 0 0.000121PF
C7_2 U237:C 0 0.000045PF
C8_2 iDFF_1_q_reg:Q 0 0.000045PF
C9_2 INP_PNN1_15 0 0.000034PF
C10_2 INP_PNN1_14 0 0.000051PF
C11_2 INP_PNN1_13 0 0.000328PF
C12_2 INP_PNN1_12 0 0.000328PF
C13_2 INP_PNN1_10 0 0.000121PF
C14_2 U246:A 0 0.000090PF
C15_2 INP_PNN1_3 0 0.000121PF
C16_2 INP_PNN1_1 0 0.000518PF
R1_2 INP_PNN1_1 INP_PNN1_2 4.408000
R2_2 INP_PNN1_1 INP_PNN1_3 4.000000
R3_2 INP_PNN1_2 INP_PNN1_4 0.304000
R4_2 INP_PNN1_2 INP_PNN1_5 4.000000
R5_2 INP_PNN1_3 U246:A 4.000000
R6_2 INP_PNN1_4 INP_PNN1_7 4.000000
R7_2 INP_PNN1_5 U237:C 4.000000
R8_2 INP_PNN1_7 INP_PNN1_9 1.824000
R9_2 U246:A INP_PNN1_10 4.000000
R10_2 INP_PNN1_9 U248:C 4.000000
R11_2 INP_PNN1_10 INP_PNN1_12 4.000000
R12_2 INP_PNN1_13 INP_PNN1_12 1.368000
R13_2 INP_PNN1_13 INP_PNN1_14 4.000000
R14_2 INP_PNN1_15 INP_PNN1_14 0.152000
R15_2 INP_PNN1_15 iDFF_1_q_reg:Q 4.000000

C1_39 U229:A 0 0.000045PF
C2_39 INP_PNN9_12 0 0.000029PF
C3_39 INP_PNN9_10 0 0.000046PF
C4_39 INP_PNN9_8 0 0.000608PF
C5_39 INP_PNN9_5 0 0.000504PF
C6_39 INP_PNN9_2 0 0.000135PF
C7_39 INP_PNN9_4 0 0.000031PF
C8_39 U249:A 0 0.000045PF
C9_39 iDFF_3_q_reg:Q 0 0.000045PF
C10_39 INP_PNN9_13 0 0.000093PF
C11_39 INP_PNN9_11 0 0.000093PF
C12_39 INP_PNN9_9 0 0.000122PF
C13_39 U198:A 0 0.000037PF
C14_39 INP_PNN9_3 0 0.000060PF
C15_39 INP_PNN9_1 0 0.000122PF
R1_39 INP_PNN9_1 INP_PNN9_2 0.760000
R2_39 INP_PNN9_1 INP_PNN9_3 4.000000
R3_39 INP_PNN9_2 INP_PNN9_4 0.110200
R4_39 INP_PNN9_2 INP_PNN9_5 4.000000
R5_39 INP_PNN9_3 U198:A 0.304000
R6_39 INP_PNN9_4 U249:A 4.000000
R7_39 INP_PNN9_5 INP_PNN9_8 5.168000
R8_39 INP_PNN9_8 INP_PNN9_9 2.128000
R9_39 INP_PNN9_8 INP_PNN9_10 4.000000
R10_39 INP_PNN9_9 INP_PNN9_11 4.000000
R11_39 INP_PNN9_10 INP_PNN9_12 0.110200
R12_39 INP_PNN9_13 INP_PNN9_11 0.912000
R13_39 INP_PNN9_12 U229:A 4.000000
R14_39 INP_PNN9_13 iDFF_3_q_reg:Q 4.000000

C1_234 U191:Z 0 0.000045PF
C2_234 n170_6 0 0.000056PF
C3_234 n170_5 0 0.000072PF
C4_234 n170_4 0 0.000292PF
C5_234 n170_3 0 0.000292PF
C6_234 n170_2 0 0.000121PF
C7_234 U190:A 0 0.000095PF
R1_234 U190:A n170_2 2.000000
R2_234 n170_2 n170_3 4.000000
R3_234 n170_3 n170_4 1.216000
R4_234 n170_4 n170_5 4.000000
R5_234 n170_5 n170_6 0.152000
R6_234 n170_6 U191:Z 4.000000

C1_267 clk_r_REG10_S2:Q 0 0.000045PF
C2_267 n45_6 0 0.000121PF
C3_267 n45_5 0 0.000138PF
C4_267 n45_4 0 0.000138PF
C5_267 n45_3 0 0.000140PF
C6_267 n45_2 0 0.000140PF
C7_267 oDFF_3_q_reg:D 0 0.000045PF
R1_267 oDFF_3_q_reg:D n45_2 4.000000
R2_267 n45_2 n45_3 1.520000
R3_267 n45_3 n45_4 4.000000
R4_267 n45_5 n45_4 1.520000
R5_267 n45_5 n45_6 4.000000
R6_267 n45_6 clk_r_REG10_S2:Q 4.000000

C1_23 iDFF_9_q_reg:Q 0 0.000045PF
C2_23 INP_PNN33_10 0 0.000298PF
C3_23 INP_PNN33_12 0 0.000282PF
C4_23 INP_PNN33_15 0 0.000650PF
C5_23 INP_PNN33_16 0 0.000650PF
C6_23 INP_PNN33_17 0 0.000105PF
C7_23 INP_PNN33_18 0 0.000123PF
C8_23 INP_PNN33_19 0 0.000125PF
C9_23 INP_PNN33_20 0 0.000090PF
C10_23 U190:C 0 0.000045PF
C11_23 clk_r_REG26_S2:D 0 0.000045PF
C12_23 INP_PNN33_4 0 0.000057PF
C13_23 INP_PNN33_2 0 0.000148PF
C14_23 INP_PNN33_5 0 0.000310PF
C15_23 INP_PNN33_8 0 0.000310PF
C16_23 U237:B 0 0.000045PF
C17_23 INP_PNN33_11 0 0.000039PF
C18_23 INP_PNN33_9 0 0.000055PF
C19_23 INP_PNN33_6 0 0.000415PF
C20_23 INP_PNN33_3 0 0.000415PF
C21_23 INP_PNN33_1 0 0.000110PF
R1_23 INP_PNN33_2 INP_PNN33_1 1.824000
R2_23 INP_PNN33_1 INP_PNN33_3 4.000000
R3_23 INP_PNN33_4 INP_PNN33_2 0.456000
R4_23 INP_PNN33_2 INP_PNN33_5 4.000000
R5_23 INP_PNN33_6 INP_PNN33_3 2.128000
R6_23 INP_PNN33_4 clk_r_REG26_S2:D 4.000000
R7_23 INP_PNN33_5 INP_PNN33_8 2.432000
R8_23 INP_PNN33_6 INP_PNN33_9 4.000000
R9_23 INP_PNN33_8 INP_PNN33_10 4.000000
R10_23 INP_PNN33_11 INP_PNN33_9 0.152000
R11_23 INP_PNN33_10 INP_PNN33_12 3.344000
R12_23 INP_PNN33_10 iDFF_9_q_reg:Q 4.000000
R13_23 INP_PNN33_11 U237:B 4.000000
R14_23 INP_PNN33_12 INP_PNN33_15 4.000000
R15_23 INP_PNN33_15 INP_PNN33_16 2.432000
R16_23 INP_PNN33_16 INP_PNN33_17 4.000000
R17_23 INP_PNN33_17 INP_PNN33_18 0.456000
R18_23 INP_PNN33_19 INP_PNN33_18 0.152000
R19_23 INP_PNN33_20 INP_PNN33_19 0.304000
R20_23 INP_PNN33_20 U190:C 4.000000

C1_25 iDFF_11_q_reg:Q 0 0.000045PF
C2_25 INP_PNN41_9 0 0.000846PF
C3_25 INP_PNN41_11 0 0.000057PF
C4_25 INP_PNN41_13 0 0.000057PF
C5_25 INP_PNN41_14 0 0.000052PF
C6_25 INP_PNN41_15 0 0.000035PF
C7_25 clk_r_REG30_S2:D 0 0.000045PF
C8_25 U196:B 0 0.000045PF
C9_25 INP_PNN41_8 0 0.000039PF
C10_25 INP_PNN41_5 0 0.000055PF
C11_25 INP_PNN41_2 0 0.001968PF
C12_25 INP_PNN41_4 0 0.000272PF
C13_25 INP_PNN41_7 0 0.000829PF
C14_25 U191:B 0 0.000045PF
C15_25 INP_PNN41_3 0 0.000121PF
C16_25 INP_PNN41_1 0 0.001714PF
R1_25 INP_PNN41_1 INP_PNN41_2 8.056000
R2_25 INP_PNN41_1 INP_PNN41_3 4.000000
R3_25 INP_PNN41_2 INP_PNN41_4 2.736000
R4_25 INP_PNN41_2 INP_PNN41_5 4.000000
R5_25 INP_PNN41_3 U191:B 4.000000
R6_25 INP_PNN41_4 INP_PNN41_7 4.000000
R7_25 INP_PNN41_5 INP_PNN41_8 0.152000
R8_25 INP_PNN41_9 INP_PNN41_7 9.272000
R9_25 INP_PNN41_8 U196:B 4.000000
R10_25 INP_PNN41_9 INP_PNN41_11 4.000000
R11_25 INP_PNN41_9 iDFF_11_q_reg:Q 4.000000
R12_25 INP_PNN41_11 INP_PNN41_13 0.304000
R13_25 INP_PNN41_13 INP_PNN41_14 4.000000
R14_25 INP_PNN41_15 INP_PNN41_14 0.152000
R15_25 INP_PNN41_15 clk_r_REG30_S2:D 4.000000

C1_62 PNN25 0 0.001944PF
C2_62 PNN25_4 0 0.001965PF
C3_62 PNN25_3 0 0.000121PF
C4_62 PNN25_2 0 0.000659PF
C5_62 iDFF_7_q_reg:D 0 0.000637PF
R1_62 iDFF_7_q_reg:D PNN25_2 6.840000
R2_62 PNN25_2 PNN25_3 4.000000
R3_62 PNN25_3 PNN25_4 4.000000
R4_62 PNN25_4 PNN25 24.015999

C1_173 U240:B 0 0.000045PF
C2_173 n109_7 0 0.000055PF
C3_173 n109_6 0 0.000071PF
C4_173 n109_5 0 0.000204PF
C5_173 n109_4 0 0.000204PF
C6_173 n109_3 0 0.000072PF
C7_173 n109_2 0 0.000056PF
C8_173 U241:Z 0 0.000045PF
R1_173 U241:Z n109_2 4.000000
R2_173 n109_3 n109_2 0.152000
R3_173 n109_3 n109_4 4.000000
R4_173 n109_5 n109_4 1.824000
R5_173 n109_5 n109_6 4.000000
R6_173 n109_6 n109_7 0.152000
R7_173 n109_7 U240:B 4.000000

C1_281 clk_r_REG0_S2:D 0 0.000087PF
C2_281 U316:A 0 0.000055PF
C3_281 U247:A 0 0.000045PF
C4_281 n58_4 0 0.000600PF
C5_281 n58_7 0 0.000572PF
C6_281 n58_10 0 0.000128PF
C7_281 n58_12 0 0.000128PF
C8_281 n58_14 0 0.000123PF
C9_281 n58_16 0 0.000123PF
C10_281 U169:D 0 0.000045PF
C11_281 n58_13 0 0.000054PF
C12_281 n58_11 0 0.000071PF
C13_281 n58_9 0 0.000741PF
C14_281 n58_5 0 0.000741PF
C15_281 n58_2 0 0.000188PF
C16_281 U178:Z 0 0.000042PF
C17_281 n58_3 0 0.000065PF
C18_281 n58_1 0 0.000160PF
R1_281 n58_2 n58_1 1.824000
R2_281 n58_1 n58_3 4.000000
R3_281 n58_4 n58_2 0.304000
R4_281 n58_2 n58_5 4.000000
R5_281 n58_3 U178:Z 0.456000
R6_281 n58_7 n58_4 5.016000
R7_281 n58_4 U247:A 4.000000
R8_281 n58_5 n58_9 1.976000
R9_281 n58_7 n58_10 4.000000
R10_281 n58_9 n58_11 4.000000
R11_281 n58_12 n58_10 0.912000
R12_281 n58_11 n58_13 0.152000
R13_281 n58_12 n58_14 4.000000
R14_281 n58_13 U169:D 4.000000
R15_281 n58_16 n58_14 0.456000
R16_281 n58_16 clk_r_REG0_S2:D 4.000000
R17_281 U316:A clk_r_REG0_S2:D 0.608000

C1_196 U172:C 0 0.000045PF
C2_196 n130_2 0 0.000214PF
C3_196 n130_4 0 0.000088PF
C4_196 n130_6 0 0.000088PF
C5_196 n130_7 0 0.000154PF
C6_196 n130_8 0 0.000201PF
C7_196 U192:Z 0 0.000095PF
C8_196 U175:C 0 0.000045PF
C9_196 n130_1 0 0.000214PF
R1_196 n130_2 n130_1 1.976000
R2_196 n130_1 U175:C 4.000000
R3_196 n130_2 n130_4 4.000000
R4_196 n130_2 U172:C 4.000000
R5_196 n130_6 n130_4 0.304000
R6_196 n130_6 n130_7 4.000000
R7_196 n130_8 n130_7 1.520000
R8_196 n130_8 U192:Z 2.000000

C1_191 U194:Z 0 0.000045PF
C2_191 n125_9 0 0.000121PF
C3_191 n125_7 0 0.001460PF
C4_191 n125_4 0 0.001460PF
C5_191 n125_2 0 0.000086PF
C6_191 U173:C 0 0.000045PF
C7_191 U171:C 0 0.000045PF
C8_191 n125_6 0 0.000146PF
C9_191 n125_3 0 0.000180PF
C10_191 n125_1 0 0.000121PF
R1_191 n125_2 n125_1 0.608000
R2_191 n125_1 n125_3 0.152000
R3_191 n125_2 n125_4 4.000000
R4_191 n125_2 U173:C 4.000000
R5_191 n125_3 n125_6 1.520000
R6_191 n125_4 n125_7 3.952000
R7_191 n125_6 U171:C 4.000000
R8_191 n125_7 n125_9 4.000000
R9_191 n125_9 U194:Z 4.000000

C1_85 U229:Z 0 0.000045PF
C2_85 Q_PNN726_5 0 0.000121PF
C3_85 Q_PNN726_4 0 0.000099PF
C4_85 Q_PNN726_3 0 0.000099PF
C5_85 Q_PNN726_2 0 0.000121PF
C6_85 clk_r_REG10_S2:D 0 0.000045PF
R1_85 clk_r_REG10_S2:D Q_PNN726_2 4.000000
R2_85 Q_PNN726_2 Q_PNN726_3 4.000000
R3_85 Q_PNN726_4 Q_PNN726_3 1.368000
R4_85 Q_PNN726_4 Q_PNN726_5 4.000000
R5_85 Q_PNN726_5 U229:Z 4.000000

C1_216 U249:Z 0 0.000045PF
C2_216 n154_8 0 0.000121PF
C3_216 n154_7 0 0.001890PF
C4_216 n154_6 0 0.001924PF
C5_216 n154_5 0 0.000393PF
C6_216 n154_4 0 0.000358PF
C7_216 n154_3 0 0.000123PF
C8_216 n154_2 0 0.000123PF
C9_216 U248:A 0 0.000045PF
R1_216 U248:A n154_2 4.000000
R2_216 n154_2 n154_3 0.456000
R3_216 n154_3 n154_4 4.000000
R4_216 n154_4 n154_5 2.280000
R5_216 n154_5 n154_6 0.152000
R6_216 n154_6 n154_7 11.248000
R7_216 n154_7 n154_8 4.000000
R8_216 n154_8 U249:Z 4.000000

C1_176 U230:Z 0 0.000079PF
C2_176 n111_6 0 0.000101PF
C3_176 n111_5 0 0.000121PF
C4_176 n111_4 0 0.000060PF
C5_176 n111_3 0 0.000060PF
C6_176 n111_2 0 0.000121PF
C7_176 U229:B 0 0.000045PF
R1_176 U229:B n111_2 4.000000
R2_176 n111_2 n111_3 4.000000
R3_176 n111_4 n111_3 0.456000
R4_176 n111_4 n111_5 4.000000
R5_176 n111_5 n111_6 4.000000
R6_176 U230:Z n111_6 0.874000

C1_187 U172:Z 0 0.000045PF
C2_187 n121_7 0 0.000052PF
C3_187 n121_6 0 0.000052PF
C4_187 n121_5 0 0.000571PF
C5_187 n121_4 0 0.000571PF
C6_187 n121_3 0 0.000194PF
C7_187 n121_2 0 0.000194PF
C8_187 U170:A 0 0.000045PF
R1_187 U170:A n121_2 4.000000
R2_187 n121_3 n121_2 1.824000
R3_187 n121_3 n121_4 4.000000
R4_187 n121_4 n121_5 2.128000
R5_187 n121_5 n121_6 4.000000
R6_187 n121_7 n121_6 0.304000
R7_187 n121_7 U172:Z 4.000000

C1_201 U196:Z 0 0.000045PF
C2_201 n139_7 0 0.000121PF
C3_201 n139_6 0 0.000155PF
C4_201 n139_5 0 0.000190PF
C5_201 n139_4 0 0.000086PF
C6_201 n139_3 0 0.000094PF
C7_201 n139_2 0 0.000094PF
C8_201 U159:C 0 0.000045PF
R1_201 U159:C n139_2 4.000000
R2_201 n139_3 n139_2 1.520000
R3_201 n139_3 n139_4 4.000000
R4_201 n139_5 n139_4 0.152000
R5_201 n139_5 n139_6 1.520000
R6_201 n139_6 n139_7 4.000000
R7_201 n139_7 U196:Z 4.000000

C1_11 U192:C 0 0.000045PF
C2_11 INP_PNN13_10 0 0.000203PF
C3_11 INP_PNN13_7 0 0.000203PF
C4_11 INP_PNN13_4 0 0.000388PF
C5_11 INP_PNN13_2 0 0.001950PF
C6_11 INP_PNN13_5 0 0.000121PF
C7_11 U248:B 0 0.000045PF
C8_11 iDFF_4_q_reg:Q 0 0.000045PF
C9_11 INP_PNN13_17 0 0.000068PF
C10_11 INP_PNN13_16 0 0.000068PF
C11_11 INP_PNN13_15 0 0.000080PF
C12_11 INP_PNN13_14 0 0.000080PF
C13_11 INP_PNN13_13 0 0.000050PF
C14_11 INP_PNN13_12 0 0.000034PF
C15_11 U240:A 0 0.000090PF
C16_11 INP_PNN13_6 0 0.000097PF
C17_11 INP_PNN13_3 0 0.000097PF
C18_11 INP_PNN13_1 0 0.001580PF
R1_11 INP_PNN13_1 INP_PNN13_2 9.728000
R2_11 INP_PNN13_1 INP_PNN13_3 4.000000
R3_11 INP_PNN13_2 INP_PNN13_4 1.824000
R4_11 INP_PNN13_2 INP_PNN13_5 4.000000
R5_11 INP_PNN13_6 INP_PNN13_3 1.064000
R6_11 INP_PNN13_4 INP_PNN13_7 4.000000
R7_11 INP_PNN13_5 U248:B 4.000000
R8_11 INP_PNN13_6 U240:A 4.000000
R9_11 INP_PNN13_10 INP_PNN13_7 2.432000
R10_11 INP_PNN13_10 U192:C 4.000000
R11_11 U240:A INP_PNN13_12 4.000000
R12_11 INP_PNN13_13 INP_PNN13_12 0.152000
R13_11 INP_PNN13_13 INP_PNN13_14 4.000000
R14_11 INP_PNN13_15 INP_PNN13_14 1.216000
R15_11 INP_PNN13_15 INP_PNN13_16 4.000000
R16_11 INP_PNN13_17 INP_PNN13_16 1.064000
R17_11 INP_PNN13_17 iDFF_4_q_reg:Q 4.000000

C1_24 U194:B 0 0.000045PF
C2_24 INP_PNN37_7 0 0.000121PF
C3_24 INP_PNN37_4 0 0.000332PF
C4_24 INP_PNN37_2 0 0.001173PF
C5_24 INP_PNN37_5 0 0.000240PF
C6_24 INP_PNN37_8 0 0.000240PF
C7_24 iDFF_10_q_reg:Q 0 0.000090PF
C8_24 INP_PNN37_11 0 0.000083PF
C9_24 INP_PNN37_12 0 0.000083PF
C10_24 INP_PNN37_13 0 0.000155PF
C11_24 INP_PNN37_14 0 0.000155PF
C12_24 INP_PNN37_15 0 0.000082PF
C13_24 INP_PNN37_16 0 0.000082PF
C14_24 clk_r_REG29_S2:D 0 0.000045PF
C15_24 U190:B 0 0.000045PF
C16_24 INP_PNN37_3 0 0.000121PF
C17_24 INP_PNN37_1 0 0.000860PF
R1_24 INP_PNN37_1 INP_PNN37_2 4.408000
R2_24 INP_PNN37_1 INP_PNN37_3 4.000000
R3_24 INP_PNN37_2 INP_PNN37_4 2.736000
R4_24 INP_PNN37_2 INP_PNN37_5 4.000000
R5_24 INP_PNN37_3 U190:B 4.000000
R6_24 INP_PNN37_4 INP_PNN37_7 4.000000
R7_24 INP_PNN37_8 INP_PNN37_5 2.128000
R8_24 INP_PNN37_7 U194:B 4.000000
R9_24 INP_PNN37_8 iDFF_10_q_reg:Q 4.000000
R10_24 iDFF_10_q_reg:Q INP_PNN37_11 4.000000
R11_24 INP_PNN37_12 INP_PNN37_11 0.760000
R12_24 INP_PNN37_12 INP_PNN37_13 4.000000
R13_24 INP_PNN37_14 INP_PNN37_13 1.064000
R14_24 INP_PNN37_14 INP_PNN37_15 4.000000
R15_24 INP_PNN37_16 INP_PNN37_15 0.912000
R16_24 INP_PNN37_16 clk_r_REG29_S2:D 4.000000

C1_186 U170:Z 0 0.000045PF
C2_186 n120_7 0 0.000149PF
C3_186 n120_6 0 0.000149PF
C4_186 n120_5 0 0.000826PF
C5_186 n120_4 0 0.000826PF
C6_186 n120_3 0 0.000245PF
C7_186 n120_2 0 0.000245PF
C8_186 U169:E 0 0.000045PF
R1_186 U169:E n120_2 4.000000
R2_186 n120_2 n120_3 0.912000
R3_186 n120_3 n120_4 4.000000
R4_186 n120_4 n120_5 3.648000
R5_186 n120_5 n120_6 4.000000
R6_186 n120_6 n120_7 1.064000
R7_186 n120_7 U170:Z 4.000000

C1_270 oDFF_4_q_reg:D 0 0.000045PF
C2_270 n48_6 0 0.000128PF
C3_270 n48_5 0 0.000128PF
C4_270 n48_4 0 0.000055PF
C5_270 n48_3 0 0.000055PF
C6_270 n48_2 0 0.000121PF
C7_270 clk_r_REG8_S2:Q 0 0.000045PF
R1_270 clk_r_REG8_S2:Q n48_2 4.000000
R2_270 n48_2 n48_3 4.000000
R3_270 n48_3 n48_4 0.608000
R4_270 n48_4 n48_5 4.000000
R5_270 n48_6 n48_5 1.824000
R6_270 n48_6 oDFF_4_q_reg:D 4.000000

C1_198 U174:Z 0 0.000045PF
C2_198 n132_6 0 0.000121PF
C3_198 n132_5 0 0.000073PF
C4_198 n132_4 0 0.000073PF
C5_198 n132_3 0 0.000199PF
C6_198 n132_2 0 0.000199PF
C7_198 U173:B 0 0.000045PF
R1_198 U173:B n132_2 4.000000
R2_198 n132_2 n132_3 1.672000
R3_198 n132_3 n132_4 4.000000
R4_198 n132_4 n132_5 0.608000
R5_198 n132_5 n132_6 4.000000
R6_198 n132_6 U174:Z 4.000000

C1_157 U175:Z 0 0.000045PF
C2_157 c0_n49_6 0 0.000054PF
C3_157 c0_n49_5 0 0.000071PF
C4_157 c0_n49_4 0 0.000864PF
C5_157 c0_n49_3 0 0.000864PF
C6_157 c0_n49_2 0 0.000121PF
C7_157 FE_OFCC0_c0_n49:A 0 0.000045PF
R1_157 FE_OFCC0_c0_n49:A c0_n49_2 4.000000
R2_157 c0_n49_2 c0_n49_3 4.000000
R3_157 c0_n49_3 c0_n49_4 4.104000
R4_157 c0_n49_4 c0_n49_5 4.000000
R5_157 c0_n49_5 c0_n49_6 0.152000
R6_157 c0_n49_6 U175:Z 4.000000

C1_200 U197:Z 0 0.000045PF
C2_200 n138_6 0 0.000121PF
C3_200 n138_5 0 0.000182PF
C4_200 n138_4 0 0.000182PF
C5_200 n138_3 0 0.000051PF
C6_200 n138_2 0 0.000035PF
C7_200 U159:B 0 0.000045PF
R1_200 U159:B n138_2 4.000000
R2_200 n138_3 n138_2 0.152000
R3_200 n138_3 n138_4 4.000000
R4_200 n138_5 n138_4 2.128000
R5_200 n138_5 n138_6 4.000000
R6_200 n138_6 U197:Z 4.000000

C1_169 U242:B 0 0.000045PF
C2_169 n105_5 0 0.000121PF
C3_169 n105_4 0 0.000242PF
C4_169 n105_3 0 0.000242PF
C5_169 n105_2 0 0.000121PF
C6_169 U243:Z 0 0.000045PF
R1_169 U243:Z n105_2 4.000000
R2_169 n105_2 n105_3 4.000000
R3_169 n105_3 n105_4 2.128000
R4_169 n105_4 n105_5 4.000000
R5_169 n105_5 U242:B 4.000000

C1_282 U185:Z 0 0.000045PF
C2_282 n59_5 0 0.000121PF
C3_282 n59_2 0 0.000974PF
C4_282 n59_4 0 0.000366PF
C5_282 n59_7 0 0.000121PF
C6_282 U165:B 0 0.000045PF
C7_282 U170:B 0 0.000045PF
C8_282 n59_6 0 0.000159PF
C9_282 n59_3 0 0.000159PF
C10_282 n59_1 0 0.000626PF
R1_282 n59_2 n59_1 6.536000
R2_282 n59_1 n59_3 4.000000
R3_282 n59_4 n59_2 1.672000
R4_282 n59_2 n59_5 4.000000
R5_282 n59_6 n59_3 0.456000
R6_282 n59_4 n59_7 4.000000
R7_282 n59_5 U185:Z 4.000000
R8_282 n59_6 U170:B 4.000000
R9_282 n59_7 U165:B 4.000000

C1_188 U171:Z 0 0.000045PF
C2_188 n122_5 0 0.000121PF
C3_188 n122_4 0 0.000915PF
C4_188 n122_3 0 0.000915PF
C5_188 n122_2 0 0.000121PF
C6_188 U170:P 0 0.000045PF
R1_188 U170:P n122_2 4.000000
R2_188 n122_2 n122_3 4.000000
R3_188 n122_3 n122_4 6.840000
R4_188 n122_4 n122_5 4.000000
R5_188 n122_5 U171:Z 4.000000

C1_89 clk_r_REG5_S2:D 0 0.000045PF
C2_89 Q_PNN730_6 0 0.000033PF
C3_89 Q_PNN730_5 0 0.000049PF
C4_89 Q_PNN730_4 0 0.000182PF
C5_89 Q_PNN730_3 0 0.000182PF
C6_89 Q_PNN730_2 0 0.000121PF
C7_89 U242:Z 0 0.000045PF
R1_89 U242:Z Q_PNN730_2 4.000000
R2_89 Q_PNN730_2 Q_PNN730_3 4.000000
R3_89 Q_PNN730_3 Q_PNN730_4 1.368000
R4_89 Q_PNN730_4 Q_PNN730_5 4.000000
R5_89 Q_PNN730_6 Q_PNN730_5 0.152000
R6_89 Q_PNN730_6 clk_r_REG5_S2:D 4.000000

C1_273 clk_r_REG5_S2:Q 0 0.000045PF
C2_273 n50_6 0 0.000121PF
C3_273 n50_5 0 0.000126PF
C4_273 n50_4 0 0.000126PF
C5_273 n50_3 0 0.000044PF
C6_273 n50_2 0 0.000044PF
C7_273 oDFF_7_q_reg:D 0 0.000045PF
R1_273 oDFF_7_q_reg:D n50_2 4.000000
R2_273 n50_2 n50_3 0.304000
R3_273 n50_3 n50_4 4.000000
R4_273 n50_5 n50_4 0.760000
R5_273 n50_5 n50_6 4.000000
R6_273 n50_6 clk_r_REG5_S2:Q 4.000000

C1_189 U171:A 0 0.000095PF
C2_189 n123_6 0 0.000121PF
C3_189 n123_5 0 0.000201PF
C4_189 n123_4 0 0.000201PF
C5_189 n123_3 0 0.000263PF
C6_189 n123_2 0 0.000263PF
C7_189 U180:Z 0 0.000045PF
R1_189 U180:Z n123_2 4.000000
R2_189 n123_3 n123_2 1.064000
R3_189 n123_3 n123_4 4.000000
R4_189 n123_5 n123_4 1.976000
R5_189 n123_5 n123_6 4.000000
R6_189 n123_6 U171:A 2.000000

C1_21 U196:C 0 0.000045PF
C2_21 INP_PNN25_8 0 0.000210PF
C3_21 INP_PNN25_5 0 0.000210PF
C4_21 INP_PNN25_2 0 0.000732PF
C5_21 INP_PNN25_4 0 0.000510PF
C6_21 INP_PNN25_7 0 0.000175PF
C7_21 INP_PNN25_9 0 0.000175PF
C8_21 U250:B 0 0.000045PF
C9_21 iDFF_7_q_reg:Q 0 0.000045PF
C10_21 INP_PNN25_16 0 0.000121PF
C11_21 INP_PNN25_15 0 0.000331PF
C12_21 INP_PNN25_14 0 0.000331PF
C13_21 INP_PNN25_13 0 0.000148PF
C14_21 INP_PNN25_11 0 0.000148PF
C15_21 U242:A 0 0.000090PF
C16_21 INP_PNN25_3 0 0.000121PF
C17_21 INP_PNN25_1 0 0.000241PF
R1_21 INP_PNN25_2 INP_PNN25_1 3.648000
R2_21 INP_PNN25_1 INP_PNN25_3 4.000000
R3_21 INP_PNN25_4 INP_PNN25_2 2.888000
R4_21 INP_PNN25_2 INP_PNN25_5 4.000000
R5_21 INP_PNN25_3 U242:A 4.000000
R6_21 INP_PNN25_4 INP_PNN25_7 4.000000
R7_21 INP_PNN25_8 INP_PNN25_5 2.432000
R8_21 INP_PNN25_7 INP_PNN25_9 1.976000
R9_21 INP_PNN25_8 U196:C 4.000000
R10_21 U242:A INP_PNN25_11 4.000000
R11_21 INP_PNN25_9 U250:B 4.000000
R12_21 INP_PNN25_13 INP_PNN25_11 1.672000
R13_21 INP_PNN25_13 INP_PNN25_14 4.000000
R14_21 INP_PNN25_14 INP_PNN25_15 3.648000
R15_21 INP_PNN25_15 INP_PNN25_16 4.000000
R16_21 INP_PNN25_16 iDFF_7_q_reg:Q 4.000000

C1_0 FE_OFCC0_c0_n49:Z 0 0.000045PF
C2_0 FE_OFCN0_c0_n49_22 0 0.000359PF
C3_0 FE_OFCN0_c0_n49_19 0 0.000359PF
C4_0 FE_OFCN0_c0_n49_14 0 0.000062PF
C5_0 FE_OFCN0_c0_n49_10 0 0.000220PF
C6_0 FE_OFCN0_c0_n49_15 0 0.000790PF
C7_0 FE_OFCN0_c0_n49_20 0 0.000790PF
C8_0 clk_r_REG23_S2:D 0 0.000045PF
C9_0 U169:B 0 0.000045PF
C10_0 FE_OFCN0_c0_n49_11 0 0.000121PF
C11_0 FE_OFCN0_c0_n49_8 0 0.001089PF
C12_0 U235:A 0 0.000045PF
C13_0 FE_OFCN0_c0_n49_28 0 0.000121PF
C14_0 FE_OFCN0_c0_n49_25 0 0.000045PF
C15_0 FE_OFCN0_c0_n49_21 0 0.000045PF
C16_0 FE_OFCN0_c0_n49_18 0 0.000336PF
C17_0 FE_OFCN0_c0_n49_13 0 0.000336PF
C18_0 U241:A 0 0.000090PF
C19_0 FE_OFCN0_c0_n49_4 0 0.000055PF
C20_0 FE_OFCN0_c0_n49_2 0 0.000197PF
C21_0 FE_OFCN0_c0_n49_5 0 0.000930PF
C22_0 U189:A 0 0.000045PF
C23_0 FE_OFCN0_c0_n49_33 0 0.000086PF
C24_0 FE_OFCN0_c0_n49_32 0 0.000086PF
C25_0 FE_OFCN0_c0_n49_31 0 0.000061PF
C26_0 FE_OFCN0_c0_n49_29 0 0.000061PF
C27_0 FE_OFCN0_c0_n49_27 0 0.000222PF
C28_0 FE_OFCN0_c0_n49_24 0 0.000222PF
C29_0 U165:A 0 0.000090PF
C30_0 FE_OFCN0_c0_n49_12 0 0.000034PF
C31_0 FE_OFCN0_c0_n49_9 0 0.000050PF
C32_0 FE_OFCN0_c0_n49_6 0 0.000042PF
C33_0 FE_OFCN0_c0_n49_3 0 0.000042PF
C34_0 FE_OFCN0_c0_n49_1 0 0.000161PF
R1_0 FE_OFCN0_c0_n49_2 FE_OFCN0_c0_n49_1 1.672000
R2_0 FE_OFCN0_c0_n49_1 FE_OFCN0_c0_n49_3 4.000000
R3_0 FE_OFCN0_c0_n49_4 FE_OFCN0_c0_n49_2 0.152000
R4_0 FE_OFCN0_c0_n49_2 FE_OFCN0_c0_n49_5 4.000000
R5_0 FE_OFCN0_c0_n49_6 FE_OFCN0_c0_n49_3 0.304000
R6_0 FE_OFCN0_c0_n49_4 U241:A 4.000000
R7_0 FE_OFCN0_c0_n49_5 FE_OFCN0_c0_n49_8 5.168000
R8_0 FE_OFCN0_c0_n49_6 FE_OFCN0_c0_n49_9 4.000000
R9_0 FE_OFCN0_c0_n49_8 FE_OFCN0_c0_n49_10 1.216000
R10_0 FE_OFCN0_c0_n49_8 FE_OFCN0_c0_n49_11 4.000000
R11_0 FE_OFCN0_c0_n49_9 FE_OFCN0_c0_n49_12 0.152000
R12_0 U241:A FE_OFCN0_c0_n49_13 4.000000
R13_0 FE_OFCN0_c0_n49_10 FE_OFCN0_c0_n49_14 0.304000
R14_0 FE_OFCN0_c0_n49_10 FE_OFCN0_c0_n49_15 4.000000
R15_0 FE_OFCN0_c0_n49_11 U169:B 4.000000
R16_0 FE_OFCN0_c0_n49_12 U165:A 4.000000
R17_0 FE_OFCN0_c0_n49_18 FE_OFCN0_c0_n49_13 3.648000
R18_0 FE_OFCN0_c0_n49_14 FE_OFCN0_c0_n49_19 4.000000
R19_0 FE_OFCN0_c0_n49_20 FE_OFCN0_c0_n49_15 5.776000
R20_0 FE_OFCN0_c0_n49_18 FE_OFCN0_c0_n49_21 4.000000
R21_0 FE_OFCN0_c0_n49_19 FE_OFCN0_c0_n49_22 1.520000
R22_0 FE_OFCN0_c0_n49_20 clk_r_REG23_S2:D 4.000000
R23_0 U165:A FE_OFCN0_c0_n49_24 4.000000
R24_0 FE_OFCN0_c0_n49_25 FE_OFCN0_c0_n49_21 0.304000
R25_0 FE_OFCN0_c0_n49_22 FE_OFCC0_c0_n49:Z 4.000000
R26_0 FE_OFCN0_c0_n49_24 FE_OFCN0_c0_n49_27 0.912000
R27_0 FE_OFCN0_c0_n49_25 FE_OFCN0_c0_n49_28 4.000000
R28_0 FE_OFCN0_c0_n49_27 FE_OFCN0_c0_n49_29 4.000000
R29_0 FE_OFCN0_c0_n49_28 U235:A 4.000000
R30_0 FE_OFCN0_c0_n49_31 FE_OFCN0_c0_n49_29 0.456000
R31_0 FE_OFCN0_c0_n49_31 FE_OFCN0_c0_n49_32 4.000000
R32_0 FE_OFCN0_c0_n49_32 FE_OFCN0_c0_n49_33 0.608000
R33_0 FE_OFCN0_c0_n49_33 U189:A 4.000000

C1_221 U251:Z 0 0.000045PF
C2_221 n159_10 0 0.000126PF
C3_221 n159_9 0 0.000126PF
C4_221 n159_8 0 0.002626PF
C5_221 n159_7 0 0.002626PF
C6_221 n159_6 0 0.000359PF
C7_221 n159_5 0 0.000359PF
C8_221 n159_4 0 0.000548PF
C9_221 n159_3 0 0.000548PF
C10_221 n159_2 0 0.000121PF
C11_221 U250:A 0 0.000045PF
R1_221 U250:A n159_2 4.000000
R2_221 n159_2 n159_3 4.000000
R3_221 n159_4 n159_3 2.432000
R4_221 n159_4 n159_5 4.000000
R5_221 n159_6 n159_5 3.800000
R6_221 n159_6 n159_7 4.000000
R7_221 n159_8 n159_7 13.376000
R8_221 n159_8 n159_9 4.000000
R9_221 n159_10 n159_9 1.216000
R10_221 n159_10 U251:Z 4.000000

C1_232 U175:B 0 0.000045PF
C2_232 n169_2 0 0.000407PF
C3_232 n169_4 0 0.000299PF
C4_232 n169_7 0 0.000123PF
C5_232 n169_9 0 0.000123PF
C6_232 n169_11 0 0.000121PF
C7_232 U172:A 0 0.000095PF
C8_232 U176:Z 0 0.000045PF
C9_232 n169_8 0 0.000121PF
C10_232 n169_6 0 0.000089PF
C11_232 n169_3 0 0.000089PF
C12_232 n169_1 0 0.000127PF
R1_232 n169_2 n169_1 1.672000
R2_232 n169_1 n169_3 4.000000
R3_232 n169_4 n169_2 2.432000
R4_232 n169_2 U175:B 4.000000
R5_232 n169_3 n169_6 0.304000
R6_232 n169_4 n169_7 4.000000
R7_232 n169_6 n169_8 4.000000
R8_232 n169_9 n169_7 0.456000
R9_232 n169_8 U176:Z 4.000000
R10_232 n169_9 n169_11 4.000000
R11_232 n169_11 U172:A 2.000000

C1_20 U244:A 0 0.000045PF
C2_20 INP_PNN21_13 0 0.000160PF
C3_20 INP_PNN21_12 0 0.000160PF
C4_20 iDFF_6_q_reg:Q 0 0.000090PF
C5_20 INP_PNN21_10 0 0.000121PF
C6_20 INP_PNN21_8 0 0.000364PF
C7_20 INP_PNN21_5 0 0.000364PF
C8_20 INP_PNN21_2 0 0.000424PF
C9_20 INP_PNN21_4 0 0.000050PF
C10_20 U250:C 0 0.000045PF
C11_20 U194:C 0 0.000045PF
C12_20 INP_PNN21_6 0 0.000097PF
C13_20 INP_PNN21_3 0 0.000101PF
C14_20 INP_PNN21_1 0 0.000397PF
R1_20 INP_PNN21_1 INP_PNN21_2 2.432000
R2_20 INP_PNN21_1 INP_PNN21_3 0.068400
R3_20 INP_PNN21_2 INP_PNN21_4 0.304000
R4_20 INP_PNN21_2 INP_PNN21_5 4.000000
R5_20 INP_PNN21_6 INP_PNN21_3 1.216000
R6_20 INP_PNN21_4 U250:C 4.000000
R7_20 INP_PNN21_5 INP_PNN21_8 3.648000
R8_20 INP_PNN21_6 U194:C 4.000000
R9_20 INP_PNN21_8 INP_PNN21_10 4.000000
R10_20 INP_PNN21_10 iDFF_6_q_reg:Q 4.000000
R11_20 iDFF_6_q_reg:Q INP_PNN21_12 4.000000
R12_20 INP_PNN21_12 INP_PNN21_13 1.672000
R13_20 INP_PNN21_13 U244:A 4.000000

C1_154 clk_r_REG3_S2:D 0 0.000045PF
C2_154 c0_n37_5 0 0.000121PF
C3_154 c0_n37_4 0 0.000222PF
C4_154 c0_n37_3 0 0.000222PF
C5_154 c0_n37_2 0 0.000121PF
C6_154 U188:Z 0 0.000045PF
R1_154 U188:Z c0_n37_2 4.000000
R2_154 c0_n37_2 c0_n37_3 4.000000
R3_154 c0_n37_4 c0_n37_3 0.912000
R4_154 c0_n37_4 c0_n37_5 4.000000
R5_154 c0_n37_5 clk_r_REG3_S2:D 4.000000

C1_197 U205:Z 0 0.000045PF
C2_197 n131_7 0 0.000186PF
C3_197 n131_6 0 0.000186PF
C4_197 n131_5 0 0.000194PF
C5_197 n131_4 0 0.000194PF
C6_197 n131_3 0 0.000061PF
C7_197 n131_2 0 0.000061PF
C8_197 U176:A 0 0.000045PF
R1_197 U176:A n131_2 4.000000
R2_197 n131_2 n131_3 0.456000
R3_197 n131_3 n131_4 4.000000
R4_197 n131_4 n131_5 1.520000
R5_197 n131_5 n131_6 4.000000
R6_197 n131_6 n131_7 1.824000
R7_197 n131_7 U205:Z 4.000000

C1_149 U189:Z 0 0.000045PF
C2_149 c0_n22_6 0 0.000121PF
C3_149 c0_n22_5 0 0.000408PF
C4_149 c0_n22_4 0 0.000408PF
C5_149 c0_n22_3 0 0.000049PF
C6_149 c0_n22_2 0 0.000032PF
C7_149 clk_r_REG21_S2:D 0 0.000045PF
R1_149 clk_r_REG21_S2:D c0_n22_2 4.000000
R2_149 c0_n22_2 c0_n22_3 0.152000
R3_149 c0_n22_3 c0_n22_4 4.000000
R4_149 c0_n22_4 c0_n22_5 3.344000
R5_149 c0_n22_5 c0_n22_6 4.000000
R6_149 c0_n22_6 U189:Z 4.000000

C1_262 clk_r_REG17_S2:Q 0 0.000045PF
C2_262 n40_6 0 0.000170PF
C3_262 n40_5 0 0.000170PF
C4_262 n40_4 0 0.000481PF
C5_262 n40_3 0 0.000481PF
C6_262 n40_2 0 0.000121PF
C7_262 U210:A 0 0.000045PF
R1_262 U210:A n40_2 4.000000
R2_262 n40_2 n40_3 4.000000
R3_262 n40_4 n40_3 3.192000
R4_262 n40_4 n40_5 4.000000
R5_262 n40_5 n40_6 1.520000
R6_262 n40_6 clk_r_REG17_S2:Q 4.000000

C1_163 U210:B 0 0.000045PF
C2_163 n10_7 0 0.000121PF
C3_163 n10_6 0 0.000286PF
C4_163 n10_4 0 0.000286PF
C5_163 n10_2 0 0.000332PF
C6_163 U211:B 0 0.000045PF
C7_163 clk_r_REG4_S2:Q 0 0.000045PF
C8_163 n10_1 0 0.000315PF
R1_163 n10_2 n10_1 3.496000
R2_163 n10_1 clk_r_REG4_S2:Q 4.000000
R3_163 n10_2 n10_4 4.000000
R4_163 n10_2 U211:B 4.000000
R5_163 n10_6 n10_4 3.496000
R6_163 n10_6 n10_7 4.000000
R7_163 n10_7 U210:B 4.000000

C1_204 U225:Z 0 0.000045PF
C2_204 n141_7 0 0.000205PF
C3_204 n141_6 0 0.000205PF
C4_204 n141_5 0 0.000146PF
C5_204 n141_4 0 0.000146PF
C6_204 n141_3 0 0.000380PF
C7_204 n141_2 0 0.000380PF
C8_204 U197:A 0 0.000045PF
R1_204 U197:A n141_2 4.000000
R2_204 n141_2 n141_3 2.128000
R3_204 n141_3 n141_4 4.000000
R4_204 n141_4 n141_5 1.064000
R5_204 n141_5 n141_6 4.000000
R6_204 n141_6 n141_7 1.520000
R7_204 n141_7 U225:Z 4.000000

C1_224 U238:Z 0 0.000045PF
C2_224 n161_7 0 0.000055PF
C3_224 n161_6 0 0.000071PF
C4_224 n161_5 0 0.000218PF
C5_224 n161_4 0 0.000218PF
C6_224 n161_3 0 0.000125PF
C7_224 n161_2 0 0.000125PF
C8_224 U236:B 0 0.000045PF
R1_224 U236:B n161_2 4.000000
R2_224 n161_2 n161_3 1.064000
R3_224 n161_3 n161_4 4.000000
R4_224 n161_4 n161_5 2.432000
R5_224 n161_5 n161_6 4.000000
R6_224 n161_6 n161_7 0.152000
R7_224 n161_7 U238:Z 4.000000

C1_14 iDFF_36_q_reg:Q 0 0.000045PF
C2_14 INP_PNN132_7 0 0.000131PF
C3_14 INP_PNN132_6 0 0.000131PF
C4_14 INP_PNN132_5 0 0.000290PF
C5_14 INP_PNN132_4 0 0.000290PF
C6_14 INP_PNN132_3 0 0.000068PF
C7_14 INP_PNN132_2 0 0.000068PF
C8_14 U205:A 0 0.000045PF
R1_14 U205:A INP_PNN132_2 4.000000
R2_14 INP_PNN132_3 INP_PNN132_2 0.304000
R3_14 INP_PNN132_3 INP_PNN132_4 4.000000
R4_14 INP_PNN132_4 INP_PNN132_5 2.736000
R5_14 INP_PNN132_5 INP_PNN132_6 4.000000
R6_14 INP_PNN132_7 INP_PNN132_6 1.216000
R7_14 INP_PNN132_7 iDFF_36_q_reg:Q 4.000000

C1_192 U206:Z 0 0.000045PF
C2_192 n126_10 0 0.000033PF
C3_192 n126_9 0 0.000050PF
C4_192 n126_8 0 0.000050PF
C5_192 n126_7 0 0.000050PF
C6_192 n126_6 0 0.000146PF
C7_192 n126_5 0 0.000146PF
C8_192 U180:A 0 0.000090PF
C9_192 n126_3 0 0.000309PF
C10_192 n126_2 0 0.000309PF
C11_192 U174:A 0 0.000045PF
R1_192 U174:A n126_2 4.000000
R2_192 n126_2 n126_3 1.976000
R3_192 n126_3 U180:A 4.000000
R4_192 U180:A n126_5 4.000000
R5_192 n126_5 n126_6 1.520000
R6_192 n126_6 n126_7 4.000000
R7_192 n126_8 n126_7 0.304000
R8_192 n126_8 n126_9 4.000000
R9_192 n126_9 n126_10 0.152000
R10_192 n126_10 U206:Z 4.000000

C1_12 U206:A 0 0.000045PF
C2_12 INP_PNN130_7 0 0.000033PF
C3_12 INP_PNN130_6 0 0.000049PF
C4_12 INP_PNN130_5 0 0.000085PF
C5_12 INP_PNN130_4 0 0.000085PF
C6_12 INP_PNN130_3 0 0.000050PF
C7_12 INP_PNN130_2 0 0.000034PF
C8_12 iDFF_34_q_reg:Q 0 0.000045PF
R1_12 iDFF_34_q_reg:Q INP_PNN130_2 4.000000
R2_12 INP_PNN130_2 INP_PNN130_3 0.152000
R3_12 INP_PNN130_3 INP_PNN130_4 4.000000
R4_12 INP_PNN130_4 INP_PNN130_5 1.368000
R5_12 INP_PNN130_5 INP_PNN130_6 4.000000
R6_12 INP_PNN130_6 INP_PNN130_7 0.152000
R7_12 INP_PNN130_7 U206:A 4.000000

C1_170 U245:Z 0 0.000045PF
C2_170 n106_5 0 0.000121PF
C3_170 n106_4 0 0.000348PF
C4_170 n106_3 0 0.000348PF
C5_170 n106_2 0 0.000121PF
C6_170 U244:B 0 0.000045PF
R1_170 U244:B n106_2 4.000000
R2_170 n106_2 n106_3 4.000000
R3_170 n106_4 n106_3 1.368000
R4_170 n106_4 n106_5 4.000000
R5_170 n106_5 U245:Z 4.000000

C1_271 clk_r_REG6_S2:Q 0 0.000045PF
C2_271 n49_6 0 0.000040PF
C3_271 n49_5 0 0.000040PF
C4_271 n49_4 0 0.000191PF
C5_271 n49_3 0 0.000191PF
C6_271 n49_2 0 0.000121PF
C7_271 oDFF_6_q_reg:D 0 0.000045PF
R1_271 oDFF_6_q_reg:D n49_2 4.000000
R2_271 n49_2 n49_3 4.000000
R3_271 n49_4 n49_3 0.760000
R4_271 n49_4 n49_5 4.000000
R5_271 n49_5 n49_6 0.304000
R6_271 n49_6 clk_r_REG6_S2:Q 4.000000

C1_13 iDFF_35_q_reg:Q 0 0.000045PF
C2_13 INP_PNN131_6 0 0.000121PF
C3_13 INP_PNN131_5 0 0.001369PF
C4_13 INP_PNN131_4 0 0.001369PF
C5_13 INP_PNN131_3 0 0.000077PF
C6_13 INP_PNN131_2 0 0.000060PF
C7_13 U225:A 0 0.000045PF
R1_13 U225:A INP_PNN131_2 4.000000
R2_13 INP_PNN131_2 INP_PNN131_3 0.152000
R3_13 INP_PNN131_3 INP_PNN131_4 4.000000
R4_13 INP_PNN131_4 INP_PNN131_5 4.560000
R5_13 INP_PNN131_5 INP_PNN131_6 4.000000
R6_13 INP_PNN131_6 iDFF_35_q_reg:Q 4.000000

C1_53 PNN131 0 0.004069PF
C2_53 PNN131_6 0 0.004124PF
C3_53 PNN131_5 0 0.000381PF
C4_53 PNN131_4 0 0.000347PF
C5_53 PNN131_3 0 0.000049PF
C6_53 PNN131_2 0 0.000033PF
C7_53 iDFF_35_q_reg:D 0 0.000045PF
R1_53 iDFF_35_q_reg:D PNN131_2 4.000000
R2_53 PNN131_2 PNN131_3 0.152000
R3_53 PNN131_3 PNN131_4 4.000000
R4_53 PNN131_4 PNN131_5 1.368000
R5_53 PNN131_6 PNN131_5 0.152000
R6_53 PNN131_6 PNN131 35.111999

C1_295 U236:Z 0 0.000045PF
C2_295 n70_8 0 0.000121PF
C3_295 n70_7 0 0.000319PF
C4_295 n70_4 0 0.000319PF
C5_295 n70_2 0 0.000189PF
C6_295 U188:B 0 0.000090PF
C7_295 n70_9 0 0.000309PF
C8_295 n70_11 0 0.000309PF
C9_295 n70_12 0 0.000053PF
C10_295 n70_13 0 0.000053PF
C11_295 n70_14 0 0.000348PF
C12_295 n70_15 0 0.000348PF
C13_295 U184:B 0 0.000045PF
C14_295 U178:A 0 0.000042PF
C15_295 n70_3 0 0.000065PF
C16_295 n70_1 0 0.000189PF
R1_295 n70_1 n70_2 1.520000
R2_295 n70_1 n70_3 4.000000
R3_295 n70_2 n70_4 4.000000
R4_295 n70_2 U188:B 4.000000
R5_295 U178:A n70_3 0.456000
R6_295 n70_4 n70_7 2.736000
R7_295 n70_7 n70_8 4.000000
R8_295 U188:B n70_9 4.000000
R9_295 n70_8 U236:Z 4.000000
R10_295 n70_9 n70_11 2.432000
R11_295 n70_11 n70_12 4.000000
R12_295 n70_13 n70_12 0.456000
R13_295 n70_13 n70_14 4.000000
R14_295 n70_14 n70_15 1.368000
R15_295 n70_15 U184:B 4.000000

C1_156 clk_r_REG17_S2:D 0 0.000110PF
C2_156 U164:Z 0 0.000045PF
C3_156 c0_n47_9 0 0.001070PF
C4_156 c0_n47_8 0 0.001070PF
C5_156 c0_n47_7 0 0.000086PF
C6_156 c0_n47_6 0 0.000196PF
C7_156 c0_n47_5 0 0.000162PF
C8_156 c0_n47_3 0 0.000046PF
C9_156 c0_n47_2 0 0.000046PF
C10_156 U161:A 0 0.000155PF
R1_156 U161:A c0_n47_2 4.000000
R2_156 c0_n47_2 c0_n47_3 0.304000
R3_156 clk_r_REG17_S2:D U161:A 1.216000
R4_156 c0_n47_3 c0_n47_5 4.000000
R5_156 c0_n47_5 c0_n47_6 0.912000
R6_156 c0_n47_6 c0_n47_7 0.152000
R7_156 c0_n47_7 c0_n47_8 4.000000
R8_156 c0_n47_8 c0_n47_9 7.144000
R9_156 c0_n47_9 U164:Z 4.000000

C1_10 iDFF_33_q_reg:Q 0 0.000045PF
C2_10 INP_PNN129_7 0 0.000038PF
C3_10 INP_PNN129_6 0 0.000055PF
C4_10 INP_PNN129_5 0 0.000187PF
C5_10 INP_PNN129_4 0 0.000187PF
C6_10 INP_PNN129_3 0 0.000209PF
C7_10 INP_PNN129_2 0 0.000209PF
C8_10 U224:A 0 0.000045PF
R1_10 U224:A INP_PNN129_2 4.000000
R2_10 INP_PNN129_3 INP_PNN129_2 1.216000
R3_10 INP_PNN129_3 INP_PNN129_4 4.000000
R4_10 INP_PNN129_4 INP_PNN129_5 0.760000
R5_10 INP_PNN129_5 INP_PNN129_6 4.000000
R6_10 INP_PNN129_7 INP_PNN129_6 0.152000
R7_10 INP_PNN129_7 iDFF_33_q_reg:Q 4.000000

C1_88 U244:Z 0 0.000045PF
C2_88 Q_PNN729_7 0 0.000033PF
C3_88 Q_PNN729_6 0 0.000049PF
C4_88 Q_PNN729_5 0 0.000871PF
C5_88 Q_PNN729_4 0 0.000871PF
C6_88 Q_PNN729_3 0 0.000039PF
C7_88 Q_PNN729_2 0 0.000039PF
C8_88 clk_r_REG6_S2:D 0 0.000045PF
R1_88 clk_r_REG6_S2:D Q_PNN729_2 4.000000
R2_88 Q_PNN729_2 Q_PNN729_3 0.304000
R3_88 Q_PNN729_3 Q_PNN729_4 4.000000
R4_88 Q_PNN729_5 Q_PNN729_4 5.320000
R5_88 Q_PNN729_5 Q_PNN729_6 4.000000
R6_88 Q_PNN729_7 Q_PNN729_6 0.152000
R7_88 Q_PNN729_7 U244:Z 4.000000

C1_227 U224:Z 0 0.000045PF
C2_227 n164_7 0 0.000192PF
C3_227 n164_6 0 0.000192PF
C4_227 n164_5 0 0.000414PF
C5_227 n164_4 0 0.000414PF
C6_227 n164_3 0 0.000123PF
C7_227 n164_2 0 0.000123PF
C8_227 U238:A 0 0.000045PF
R1_227 U238:A n164_2 4.000000
R2_227 n164_2 n164_3 1.216000
R3_227 n164_3 n164_4 4.000000
R4_227 n164_4 n164_5 2.128000
R5_227 n164_5 n164_6 4.000000
R6_227 n164_6 n164_7 0.760000
R7_227 n164_7 U224:Z 4.000000

C1_250 clk_r_REG37_S2:Q 0 0.000045PF
C2_250 n29_6 0 0.000032PF
C3_250 n29_5 0 0.000049PF
C4_250 n29_4 0 0.000185PF
C5_250 n29_3 0 0.000185PF
C6_250 n29_2 0 0.000121PF
C7_250 U288:A 0 0.000045PF
R1_250 U288:A n29_2 4.000000
R2_250 n29_2 n29_3 4.000000
R3_250 n29_4 n29_3 1.368000
R4_250 n29_4 n29_5 4.000000
R5_250 n29_5 n29_6 0.152000
R6_250 n29_6 clk_r_REG37_S2:Q 4.000000

C1_150 U184:Z 0 0.000045PF
C2_150 c0_n23_6 0 0.000054PF
C3_150 c0_n23_5 0 0.000071PF
C4_150 c0_n23_4 0 0.000588PF
C5_150 c0_n23_3 0 0.000588PF
C6_150 c0_n23_2 0 0.000121PF
C7_150 clk_r_REG11_S2:D 0 0.000045PF
R1_150 clk_r_REG11_S2:D c0_n23_2 4.000000
R2_150 c0_n23_2 c0_n23_3 4.000000
R3_150 c0_n23_3 c0_n23_4 5.320000
R4_150 c0_n23_4 c0_n23_5 4.000000
R5_150 c0_n23_6 c0_n23_5 0.152000
R6_150 c0_n23_6 U184:Z 4.000000

C1_292 U308:Z 0 0.000045PF
C2_292 n68_7 0 0.000121PF
C3_292 n68_4 0 0.000150PF
C4_292 n68_2 0 0.000356PF
C5_292 n68_5 0 0.000379PF
C6_292 n68_8 0 0.000379PF
C7_292 U201:A 0 0.000045PF
C8_292 U202:A 0 0.000045PF
C9_292 n68_3 0 0.000121PF
C10_292 n68_1 0 0.000224PF
R1_292 n68_1 n68_2 0.912000
R2_292 n68_1 n68_3 4.000000
R3_292 n68_2 n68_4 0.608000
R4_292 n68_2 n68_5 4.000000
R5_292 n68_3 U202:A 4.000000
R6_292 n68_4 n68_7 4.000000
R7_292 n68_5 n68_8 3.648000
R8_292 n68_7 U308:Z 4.000000
R9_292 n68_8 U201:A 4.000000

C1_159 U183:Z 0 0.000045PF
C2_159 c0_n56_7 0 0.000232PF
C3_159 c0_n56_6 0 0.000232PF
C4_159 c0_n56_5 0 0.000353PF
C5_159 c0_n56_4 0 0.000353PF
C6_159 c0_n56_3 0 0.000051PF
C7_159 c0_n56_2 0 0.000035PF
C8_159 clk_r_REG4_S2:D 0 0.000045PF
R1_159 clk_r_REG4_S2:D c0_n56_2 4.000000
R2_159 c0_n56_2 c0_n56_3 0.152000
R3_159 c0_n56_3 c0_n56_4 4.000000
R4_159 c0_n56_4 c0_n56_5 1.520000
R5_159 c0_n56_5 c0_n56_6 4.000000
R6_159 c0_n56_6 c0_n56_7 1.824000
R7_159 c0_n56_7 U183:Z 4.000000

C1_19 U226:B 0 0.000045PF
C2_19 INP_PNN137_14 0 0.000121PF
C3_19 INP_PNN137_9 0 0.000125PF
C4_19 INP_PNN137_7 0 0.000214PF
C5_19 INP_PNN137_10 0 0.000128PF
C6_19 INP_PNN137_15 0 0.000128PF
C7_19 U206:B 0 0.000045PF
C8_19 iDFF_41_q_reg:Q 0 0.000045PF
C9_19 INP_PNN137_24 0 0.000220PF
C10_19 INP_PNN137_18 0 0.000075PF
C11_19 INP_PNN137_13 0 0.000642PF
C12_19 U225:B 0 0.000045PF
C13_19 INP_PNN137_34 0 0.000039PF
C14_19 INP_PNN137_33 0 0.000055PF
C15_19 INP_PNN137_32 0 0.000399PF
C16_19 INP_PNN137_31 0 0.000399PF
C17_19 INP_PNN137_27 0 0.000164PF
C18_19 U227:B 0 0.000045PF
C19_19 INP_PNN137_26 0 0.000192PF
C20_19 INP_PNN137_23 0 0.000192PF
C21_19 INP_PNN137_17 0 0.000580PF
C22_19 U205:B 0 0.000045PF
C23_19 INP_PNN137_16 0 0.000170PF
C24_19 INP_PNN137_12 0 0.000170PF
C25_19 INP_PNN137_8 0 0.000407PF
C26_19 INP_PNN137_6 0 0.000291PF
C27_19 INP_PNN137_4 0 0.000050PF
C28_19 INP_PNN137_2 0 0.000218PF
C29_19 INP_PNN137_5 0 0.000171PF
C30_19 U231:A 0 0.000045PF
C31_19 INP_PNN137_25 0 0.000179PF
C32_19 INP_PNN137_21 0 0.000179PF
C33_19 U224:B 0 0.000158PF
C34_19 U228:B 0 0.000045PF
C35_19 INP_PNN137_1 0 0.000187PF
R1_19 INP_PNN137_2 INP_PNN137_1 1.824000
R2_19 INP_PNN137_1 U228:B 4.000000
R3_19 INP_PNN137_4 INP_PNN137_2 0.304000
R4_19 INP_PNN137_2 INP_PNN137_5 4.000000
R5_19 INP_PNN137_4 INP_PNN137_6 4.000000
R6_19 INP_PNN137_5 INP_PNN137_7 1.976000
R7_19 INP_PNN137_8 INP_PNN137_6 2.888000
R8_19 INP_PNN137_7 INP_PNN137_9 0.760000
R9_19 INP_PNN137_7 INP_PNN137_10 4.000000
R10_19 U224:B INP_PNN137_8 1.216000
R11_19 INP_PNN137_8 INP_PNN137_12 4.000000
R12_19 INP_PNN137_9 INP_PNN137_13 0.760000
R13_19 INP_PNN137_9 INP_PNN137_14 4.000000
R14_19 INP_PNN137_15 INP_PNN137_10 1.824000
R15_19 INP_PNN137_16 INP_PNN137_12 1.520000
R16_19 INP_PNN137_13 INP_PNN137_17 3.800000
R17_19 INP_PNN137_13 INP_PNN137_18 4.000000
R18_19 INP_PNN137_14 U226:B 4.000000
R19_19 INP_PNN137_15 U206:B 4.000000
R20_19 U224:B INP_PNN137_21 4.000000
R21_19 INP_PNN137_16 U205:B 4.000000
R22_19 INP_PNN137_17 INP_PNN137_23 4.000000
R23_19 INP_PNN137_24 INP_PNN137_18 0.456000
R24_19 INP_PNN137_21 INP_PNN137_25 1.824000
R25_19 INP_PNN137_23 INP_PNN137_26 1.824000
R26_19 INP_PNN137_27 INP_PNN137_24 1.216000
R27_19 INP_PNN137_24 iDFF_41_q_reg:Q 4.000000
R28_19 INP_PNN137_25 U231:A 4.000000
R29_19 INP_PNN137_26 U227:B 4.000000
R30_19 INP_PNN137_27 INP_PNN137_31 4.000000
R31_19 INP_PNN137_31 INP_PNN137_32 1.520000
R32_19 INP_PNN137_32 INP_PNN137_33 4.000000
R33_19 INP_PNN137_34 INP_PNN137_33 0.152000
R34_19 INP_PNN137_34 U225:B 4.000000

C1_293 U169:Z 0 0.000045PF
C2_293 n69_9 0 0.000244PF
C3_293 n69_7 0 0.000278PF
C4_293 n69_4 0 0.000886PF
C5_293 n69_2 0 0.000893PF
C6_293 U162:B 0 0.000045PF
C7_293 U183:B 0 0.000045PF
C8_293 n69_10 0 0.000437PF
C9_293 n69_8 0 0.000437PF
C10_293 n69_6 0 0.000415PF
C11_293 n69_3 0 0.000415PF
C12_293 n69_1 0 0.000060PF
R1_293 n69_2 n69_1 0.304000
R2_293 n69_1 n69_3 4.000000
R3_293 n69_4 n69_2 5.776000
R4_293 n69_2 U162:B 4.000000
R5_293 n69_3 n69_6 2.736000
R6_293 n69_4 n69_7 0.152000
R7_293 n69_6 n69_8 4.000000
R8_293 n69_9 n69_7 1.672000
R9_293 n69_8 n69_10 1.824000
R10_293 n69_9 U169:Z 4.000000
R11_293 n69_10 U183:B 4.000000

C1_318 U289:Z 0 0.000045PF
C2_318 n91_7 0 0.000148PF
C3_318 n91_6 0 0.000148PF
C4_318 n91_5 0 0.000089PF
C5_318 n91_4 0 0.000089PF
C6_318 n91_3 0 0.000050PF
C7_318 n91_2 0 0.000033PF
C8_318 U288:B 0 0.000045PF
R1_318 U288:B n91_2 4.000000
R2_318 n91_2 n91_3 0.152000
R3_318 n91_3 n91_4 4.000000
R4_318 n91_5 n91_4 0.304000
R5_318 n91_5 n91_6 4.000000
R6_318 n91_6 n91_7 1.672000
R7_318 n91_7 U289:Z 4.000000

C1_100 oDFF_18_q_reg:D 0 0.000045PF
C2_100 Q_PNN741_6 0 0.000045PF
C3_100 Q_PNN741_5 0 0.000045PF
C4_100 Q_PNN741_4 0 0.000193PF
C5_100 Q_PNN741_3 0 0.000193PF
C6_100 Q_PNN741_2 0 0.000121PF
C7_100 U288:Z 0 0.000045PF
R1_100 U288:Z Q_PNN741_2 4.000000
R2_100 Q_PNN741_2 Q_PNN741_3 4.000000
R3_100 Q_PNN741_3 Q_PNN741_4 0.912000
R4_100 Q_PNN741_4 Q_PNN741_5 4.000000
R5_100 Q_PNN741_6 Q_PNN741_5 0.304000
R6_100 Q_PNN741_6 oDFF_18_q_reg:D 4.000000

C1_104 U280:Z 0 0.000045PF
C2_104 Q_PNN745_7 0 0.000032PF
C3_104 Q_PNN745_6 0 0.000049PF
C4_104 Q_PNN745_5 0 0.000100PF
C5_104 Q_PNN745_4 0 0.000100PF
C6_104 Q_PNN745_3 0 0.000149PF
C7_104 Q_PNN745_2 0 0.000149PF
C8_104 oDFF_22_q_reg:D 0 0.000045PF
R1_104 oDFF_22_q_reg:D Q_PNN745_2 4.000000
R2_104 Q_PNN745_2 Q_PNN745_3 1.672000
R3_104 Q_PNN745_3 Q_PNN745_4 4.000000
R4_104 Q_PNN745_4 Q_PNN745_5 1.064000
R5_104 Q_PNN745_5 Q_PNN745_6 4.000000
R6_104 Q_PNN745_6 Q_PNN745_7 0.152000
R7_104 Q_PNN745_7 U280:Z 4.000000

C1_316 U203:A 0 0.000045PF
C2_316 n9_8 0 0.000039PF
C3_316 n9_5 0 0.000056PF
C4_316 n9_2 0 0.000278PF
C5_316 n9_4 0 0.000110PF
C6_316 n9_7 0 0.000056PF
C7_316 n9_10 0 0.000039PF
C8_316 U204:A 0 0.000045PF
C9_316 clk_r_REG11_S2:Q 0 0.000045PF
C10_316 n9_6 0 0.000129PF
C11_316 n9_3 0 0.000129PF
C12_316 n9_1 0 0.000187PF
R1_316 n9_1 n9_2 1.824000
R2_316 n9_1 n9_3 4.000000
R3_316 n9_2 n9_4 0.760000
R4_316 n9_2 n9_5 4.000000
R5_316 n9_6 n9_3 1.368000
R6_316 n9_4 n9_7 4.000000
R7_316 n9_5 n9_8 0.152000
R8_316 n9_6 clk_r_REG11_S2:Q 4.000000
R9_316 n9_7 n9_10 0.152000
R10_316 n9_8 U203:A 4.000000
R11_316 n9_10 U204:A 4.000000

C1_291 U204:B 0 0.000045PF
C2_291 n67_10 0 0.000039PF
C3_291 n67_9 0 0.000055PF
C4_291 n67_8 0 0.000164PF
C5_291 n67_7 0 0.000164PF
C6_291 n67_6 0 0.000219PF
C7_291 n67_4 0 0.000219PF
C8_291 U314:Z 0 0.000045PF
C9_291 n67_3 0 0.000126PF
C10_291 n67_2 0 0.000126PF
C11_291 U202:B 0 0.000090PF
R1_291 U202:B n67_2 4.000000
R2_291 n67_3 n67_2 1.216000
R3_291 U202:B n67_4 4.000000
R4_291 n67_3 U314:Z 4.000000
R5_291 n67_4 n67_6 1.824000
R6_291 n67_6 n67_7 4.000000
R7_291 n67_8 n67_7 1.216000
R8_291 n67_8 n67_9 4.000000
R9_291 n67_9 n67_10 0.152000
R10_291 n67_10 U204:B 4.000000

C1_184 U190:Z 0 0.000045PF
C2_184 n119_12 0 0.000450PF
C3_184 n119_11 0 0.000450PF
C4_184 n119_10 0 0.000057PF
C5_184 n119_9 0 0.000057PF
C6_184 n119_8 0 0.000375PF
C7_184 n119_7 0 0.000375PF
C8_184 U218:B 0 0.000090PF
C9_184 n119_5 0 0.000121PF
C10_184 n119_4 0 0.000326PF
C11_184 n119_3 0 0.000326PF
C12_184 n119_2 0 0.000121PF
C13_184 U258:B 0 0.000045PF
R1_184 U258:B n119_2 4.000000
R2_184 n119_2 n119_3 4.000000
R3_184 n119_4 n119_3 1.368000
R4_184 n119_4 n119_5 4.000000
R5_184 n119_5 U218:B 4.000000
R6_184 U218:B n119_7 4.000000
R7_184 n119_8 n119_7 4.104000
R8_184 n119_8 n119_9 4.000000
R9_184 n119_10 n119_9 0.304000
R10_184 n119_10 n119_11 4.000000
R11_184 n119_12 n119_11 5.776000
R12_184 n119_12 U190:Z 4.000000

C1_16 iDFF_38_q_reg:Q 0 0.000045PF
C2_16 INP_PNN134_6 0 0.000136PF
C3_16 INP_PNN134_5 0 0.000136PF
C4_16 INP_PNN134_4 0 0.000379PF
C5_16 INP_PNN134_3 0 0.000379PF
C6_16 INP_PNN134_2 0 0.000121PF
C7_16 U228:A 0 0.000045PF
R1_16 U228:A INP_PNN134_2 4.000000
R2_16 INP_PNN134_2 INP_PNN134_3 4.000000
R3_16 INP_PNN134_3 INP_PNN134_4 1.976000
R4_16 INP_PNN134_4 INP_PNN134_5 4.000000
R5_16 INP_PNN134_6 INP_PNN134_5 1.520000
R6_16 INP_PNN134_6 iDFF_38_q_reg:Q 4.000000

C1_312 U281:Z 0 0.000045PF
C2_312 n86_5 0 0.000121PF
C3_312 n86_4 0 0.000166PF
C4_312 n86_3 0 0.000166PF
C5_312 n86_2 0 0.000121PF
C6_312 U280:B 0 0.000045PF
R1_312 U280:B n86_2 4.000000
R2_312 n86_2 n86_3 4.000000
R3_312 n86_4 n86_3 2.128000
R4_312 n86_4 n86_5 4.000000
R5_312 n86_5 U281:Z 4.000000

C1_210 U248:Z 0 0.000045PF
C2_210 n148_12 0 0.001031PF
C3_210 n148_10 0 0.001031PF
C4_210 n148_8 0 0.000307PF
C5_210 n148_6 0 0.000307PF
C6_210 n148_4 0 0.000053PF
C7_210 n148_2 0 0.000122PF
C8_210 n148_5 0 0.001158PF
C9_210 n148_7 0 0.001158PF
C10_210 n148_9 0 0.000121PF
C11_210 U222:B 0 0.000045PF
C12_210 U216:A 0 0.000045PF
C13_210 n148_1 0 0.000088PF
R1_210 n148_2 n148_1 1.520000
R2_210 n148_1 U216:A 4.000000
R3_210 n148_4 n148_2 0.456000
R4_210 n148_2 n148_5 4.000000
R5_210 n148_4 n148_6 4.000000
R6_210 n148_5 n148_7 7.600000
R7_210 n148_8 n148_6 3.192000
R8_210 n148_7 n148_9 4.000000
R9_210 n148_8 n148_10 4.000000
R10_210 n148_9 U222:B 4.000000
R11_210 n148_12 n148_10 9.576000
R12_210 n148_12 U248:Z 4.000000

C1_17 iDFF_39_q_reg:Q 0 0.000045PF
C2_17 INP_PNN135_6 0 0.000034PF
C3_17 INP_PNN135_5 0 0.000050PF
C4_17 INP_PNN135_4 0 0.000197PF
C5_17 INP_PNN135_3 0 0.000197PF
C6_17 INP_PNN135_2 0 0.000121PF
C7_17 U231:B 0 0.000045PF
R1_17 U231:B INP_PNN135_2 4.000000
R2_17 INP_PNN135_2 INP_PNN135_3 4.000000
R3_17 INP_PNN135_4 INP_PNN135_3 0.760000
R4_17 INP_PNN135_4 INP_PNN135_5 4.000000
R5_17 INP_PNN135_5 INP_PNN135_6 0.152000
R6_17 INP_PNN135_6 iDFF_39_q_reg:Q 4.000000

C1_278 clk_r_REG28_S2:Q 0 0.000045PF
C2_278 n55_6 0 0.000032PF
C3_278 n55_5 0 0.000049PF
C4_278 n55_4 0 0.000239PF
C5_278 n55_3 0 0.000239PF
C6_278 n55_2 0 0.000121PF
C7_278 U311:A 0 0.000045PF
R1_278 U311:A n55_2 4.000000
R2_278 n55_2 n55_3 4.000000
R3_278 n55_4 n55_3 1.976000
R4_278 n55_4 n55_5 4.000000
R5_278 n55_5 n55_6 0.152000
R6_278 n55_6 clk_r_REG28_S2:Q 4.000000

C1_261 U202:C 0 0.000045PF
C2_261 n4_9 0 0.000200PF
C3_261 n4_8 0 0.000200PF
C4_261 clk_r_REG14_S2:Q 0 0.000090PF
C5_261 n4_6 0 0.000121PF
C6_261 n4_5 0 0.000111PF
C7_261 n4_4 0 0.000111PF
C8_261 n4_3 0 0.000155PF
C9_261 n4_2 0 0.000155PF
C10_261 U201:C 0 0.000045PF
R1_261 U201:C n4_2 4.000000
R2_261 n4_3 n4_2 1.368000
R3_261 n4_3 n4_4 4.000000
R4_261 n4_5 n4_4 0.760000
R5_261 n4_5 n4_6 4.000000
R6_261 n4_6 clk_r_REG14_S2:Q 4.000000
R7_261 clk_r_REG14_S2:Q n4_8 4.000000
R8_261 n4_9 n4_8 1.520000
R9_261 n4_9 U202:C 4.000000

C1_280 clk_r_REG12_S2:D 0 0.000045PF
C2_280 n57_9 0 0.000419PF
C3_280 n57_8 0 0.000419PF
C4_280 n57_7 0 0.000513PF
C5_280 n57_6 0 0.000513PF
C6_280 n57_5 0 0.000121PF
C7_280 U187:Z 0 0.000090PF
C8_280 n57_3 0 0.000252PF
C9_280 n57_2 0 0.000252PF
C10_280 U162:A 0 0.000045PF
R1_280 U162:A n57_2 4.000000
R2_280 n57_2 n57_3 1.824000
R3_280 n57_3 U187:Z 4.000000
R4_280 U187:Z n57_5 4.000000
R5_280 n57_5 n57_6 4.000000
R6_280 n57_7 n57_6 3.800000
R7_280 n57_7 n57_8 4.000000
R8_280 n57_8 n57_9 5.320000
R9_280 n57_9 clk_r_REG12_S2:D 4.000000

C1_206 U222:Z 0 0.000045PF
C2_206 n144_6 0 0.000121PF
C3_206 n144_5 0 0.000050PF
C4_206 n144_4 0 0.000050PF
C5_206 n144_3 0 0.000143PF
C6_206 n144_2 0 0.000143PF
C7_206 U220:B 0 0.000045PF
R1_206 U220:B n144_2 4.000000
R2_206 n144_3 n144_2 2.128000
R3_206 n144_3 n144_4 4.000000
R4_206 n144_5 n144_4 0.304000
R5_206 n144_5 n144_6 4.000000
R6_206 n144_6 U222:Z 4.000000

C1_144 oDFF_30_q_reg:Q 0 0.000045PF
C2_144 Qout_PNN753_4 0 0.000033PF
C3_144 Qout_PNN753_3 0 0.000049PF
C4_144 Qout_PNN753_2 0 0.003308PF
C5_144 Qout_PNN753 0 0.003287PF
R1_144 Qout_PNN753 Qout_PNN753_2 30.551999
R2_144 Qout_PNN753_2 Qout_PNN753_3 4.000000
R3_144 Qout_PNN753_4 Qout_PNN753_3 0.152000
R4_144 Qout_PNN753_4 oDFF_30_q_reg:Q 4.000000

C1_215 U218:A 0 0.000045PF
C2_215 n152_5 0 0.000121PF
C3_215 n152_4 0 0.000163PF
C4_215 n152_3 0 0.000163PF
C5_215 n152_2 0 0.000121PF
C6_215 U231:Z 0 0.000045PF
R1_215 U231:Z n152_2 4.000000
R2_215 n152_2 n152_3 4.000000
R3_215 n152_3 n152_4 1.064000
R4_215 n152_4 n152_5 4.000000
R5_215 n152_5 U218:A 4.000000

C1_286 U311:Z 0 0.000045PF
C2_286 n62_5 0 0.000121PF
C3_286 n62_2 0 0.000285PF
C4_286 n62_4 0 0.000134PF
C5_286 n62_7 0 0.000105PF
C6_286 n62_9 0 0.000070PF
C7_286 n62_10 0 0.000121PF
C8_286 U281:B 0 0.000045PF
C9_286 U289:A 0 0.000045PF
C10_286 n62_3 0 0.000121PF
C11_286 n62_1 0 0.000204PF
R1_286 n62_1 n62_2 0.912000
R2_286 n62_1 n62_3 4.000000
R3_286 n62_2 n62_4 1.216000
R4_286 n62_2 n62_5 4.000000
R5_286 n62_3 U289:A 4.000000
R6_286 n62_4 n62_7 0.152000
R7_286 n62_5 U311:Z 4.000000
R8_286 n62_7 n62_9 0.608000
R9_286 n62_9 n62_10 4.000000
R10_286 n62_10 U281:B 4.000000

C1_155 U186:Z 0 0.000045PF
C2_155 c0_n46_8 0 0.000091PF
C3_155 c0_n46_7 0 0.000091PF
C4_155 c0_n46_6 0 0.000094PF
C5_155 c0_n46_5 0 0.000094PF
C6_155 c0_n46_4 0 0.000411PF
C7_155 c0_n46_3 0 0.000411PF
C8_155 U163:A 0 0.000103PF
C9_155 clk_r_REG18_S2:D 0 0.000071PF
R1_155 U163:A clk_r_REG18_S2:D 0.760000
R2_155 U163:A c0_n46_3 4.000000
R3_155 c0_n46_3 c0_n46_4 4.560000
R4_155 c0_n46_4 c0_n46_5 4.000000
R5_155 c0_n46_6 c0_n46_5 0.760000
R6_155 c0_n46_6 c0_n46_7 4.000000
R7_155 c0_n46_7 c0_n46_8 0.608000
R8_155 c0_n46_8 U186:Z 4.000000

C1_194 U172:B 0 0.000045PF
C2_194 n129_18 0 0.000121PF
C3_194 n129_17 0 0.000239PF
C4_194 n129_16 0 0.000239PF
C5_194 n129_14 0 0.000201PF
C6_194 n129_13 0 0.000301PF
C7_194 U175:A 0 0.000045PF
C8_194 U238:B 0 0.000045PF
C9_194 n129_2 0 0.000636PF
C10_194 n129_4 0 0.000277PF
C11_194 n129_7 0 0.000496PF
C12_194 n129_9 0 0.000496PF
C13_194 n129_11 0 0.000118PF
C14_194 U212:Z 0 0.000045PF
C15_194 n129_10 0 0.000237PF
C16_194 n129_8 0 0.000237PF
C17_194 n129_6 0 0.000997PF
C18_194 n129_3 0 0.000997PF
C19_194 n129_1 0 0.000378PF
R1_194 n129_2 n129_1 4.712000
R2_194 n129_1 n129_3 4.000000
R3_194 n129_4 n129_2 2.736000
R4_194 n129_2 U238:B 4.000000
R5_194 n129_3 n129_6 10.640000
R6_194 n129_4 n129_7 4.000000
R7_194 n129_6 n129_8 4.000000
R8_194 n129_7 n129_9 2.128000
R9_194 n129_8 n129_10 3.192000
R10_194 n129_9 n129_11 4.000000
R11_194 n129_10 U212:Z 4.000000
R12_194 n129_13 n129_11 1.216000
R13_194 n129_14 n129_13 1.520000
R14_194 n129_13 U175:A 4.000000
R15_194 n129_14 n129_16 4.000000
R16_194 n129_17 n129_16 0.912000
R17_194 n129_17 n129_18 4.000000
R18_194 n129_18 U172:B 4.000000

C1_220 U227:Z 0 0.000045PF
C2_220 n158_7 0 0.000122PF
C3_220 n158_6 0 0.000122PF
C4_220 n158_5 0 0.000992PF
C5_220 n158_4 0 0.000992PF
C6_220 n158_3 0 0.000100PF
C7_220 n158_2 0 0.000100PF
C8_220 U208:A 0 0.000045PF
R1_220 U208:A n158_2 4.000000
R2_220 n158_3 n158_2 1.216000
R3_220 n158_3 n158_4 4.000000
R4_220 n158_4 n158_5 6.080000
R5_220 n158_5 n158_6 4.000000
R6_220 n158_7 n158_6 0.760000
R7_220 n158_7 U227:Z 4.000000

C1_18 iDFF_40_q_reg:Q 0 0.000045PF
C2_18 INP_PNN136_7 0 0.000046PF
C3_18 INP_PNN136_6 0 0.000046PF
C4_18 INP_PNN136_5 0 0.000561PF
C5_18 INP_PNN136_4 0 0.000561PF
C6_18 INP_PNN136_3 0 0.000143PF
C7_18 INP_PNN136_2 0 0.000143PF
C8_18 U227:A 0 0.000045PF
R1_18 U227:A INP_PNN136_2 4.000000
R2_18 INP_PNN136_2 INP_PNN136_3 1.064000
R3_18 INP_PNN136_3 INP_PNN136_4 4.000000
R4_18 INP_PNN136_4 INP_PNN136_5 2.432000
R5_18 INP_PNN136_5 INP_PNN136_6 4.000000
R6_18 INP_PNN136_6 INP_PNN136_7 0.304000
R7_18 INP_PNN136_7 iDFF_40_q_reg:Q 4.000000

C1_152 clk_r_REG14_S2:D 0 0.000110PF
C2_152 c0_n30_5 0 0.000132PF
C3_152 c0_n30_2 0 0.000371PF
C4_152 c0_n30_4 0 0.000205PF
C5_152 U184:A 0 0.000045PF
C6_152 U166:Z 0 0.000045PF
C7_152 c0_n30_10 0 0.000038PF
C8_152 c0_n30_9 0 0.000055PF
C9_152 c0_n30_6 0 0.000411PF
C10_152 c0_n30_3 0 0.000411PF
C11_152 c0_n30_1 0 0.000185PF
R1_152 c0_n30_2 c0_n30_1 1.368000
R2_152 c0_n30_1 c0_n30_3 4.000000
R3_152 c0_n30_4 c0_n30_2 1.824000
R4_152 c0_n30_2 c0_n30_5 4.000000
R5_152 c0_n30_3 c0_n30_6 4.560000
R6_152 c0_n30_4 U184:A 4.000000
R7_152 clk_r_REG14_S2:D c0_n30_5 1.216000
R8_152 c0_n30_6 c0_n30_9 4.000000
R9_152 c0_n30_9 c0_n30_10 0.152000
R10_152 c0_n30_10 U166:Z 4.000000

C1_179 U256:A 0 0.000095PF
C2_179 n114_10 0 0.000121PF
C3_179 n114_8 0 0.000155PF
C4_179 n114_6 0 0.000155PF
C5_179 n114_4 0 0.000121PF
C6_179 U252:Z 0 0.000045PF
C7_179 n114_11 0 0.000196PF
C8_179 n114_9 0 0.000230PF
C9_179 n114_7 0 0.000337PF
C10_179 n114_5 0 0.000337PF
C11_179 n114_3 0 0.001197PF
C12_179 n114_2 0 0.001162PF
C13_179 U160:A 0 0.000090PF
R1_179 U160:A n114_2 4.000000
R2_179 n114_3 n114_2 9.576000
R3_179 U160:A n114_4 4.000000
R4_179 n114_5 n114_3 0.152000
R5_179 n114_4 n114_6 4.000000
R6_179 n114_7 n114_5 2.888000
R7_179 n114_8 n114_6 1.064000
R8_179 n114_9 n114_7 0.152000
R9_179 n114_8 n114_10 4.000000
R10_179 n114_11 n114_9 2.888000
R11_179 n114_10 U256:A 2.000000
R12_179 n114_11 U252:Z 4.000000

C1_37 clk_r_REG41_S2:D 0 0.000045PF
C2_37 INP_PNN85_8 0 0.000060PF
C3_37 INP_PNN85_5 0 0.000060PF
C4_37 INP_PNN85_2 0 0.001621PF
C5_37 INP_PNN85_4 0 0.001540PF
C6_37 INP_PNN85_7 0 0.000121PF
C7_37 U259:A 0 0.000090PF
C8_37 INP_PNN85_14 0 0.000329PF
C9_37 INP_PNN85_15 0 0.000329PF
C10_37 U212:B 0 0.000045PF
C11_37 iDFF_22_q_reg:Q 0 0.000045PF
C12_37 INP_PNN85_12 0 0.000041PF
C13_37 INP_PNN85_9 0 0.000041PF
C14_37 INP_PNN85_6 0 0.000203PF
C15_37 INP_PNN85_3 0 0.000237PF
C16_37 INP_PNN85_1 0 0.000134PF
R1_37 INP_PNN85_2 INP_PNN85_1 1.672000
R2_37 INP_PNN85_3 INP_PNN85_1 0.152000
R3_37 INP_PNN85_4 INP_PNN85_2 8.208000
R4_37 INP_PNN85_2 INP_PNN85_5 4.000000
R5_37 INP_PNN85_3 INP_PNN85_6 1.064000
R6_37 INP_PNN85_4 INP_PNN85_7 4.000000
R7_37 INP_PNN85_5 INP_PNN85_8 0.456000
R8_37 INP_PNN85_6 INP_PNN85_9 4.000000
R9_37 INP_PNN85_7 U259:A 4.000000
R10_37 INP_PNN85_8 clk_r_REG41_S2:D 4.000000
R11_37 INP_PNN85_9 INP_PNN85_12 0.304000
R12_37 INP_PNN85_12 iDFF_22_q_reg:Q 4.000000
R13_37 U259:A INP_PNN85_14 4.000000
R14_37 INP_PNN85_14 INP_PNN85_15 1.520000
R15_37 INP_PNN85_15 U212:B 4.000000

C1_246 clk_r_REG41_S2:Q 0 0.000045PF
C2_246 n25_7 0 0.000034PF
C3_246 n25_6 0 0.000050PF
C4_246 n25_5 0 0.000287PF
C5_246 n25_4 0 0.000287PF
C6_246 n25_3 0 0.000092PF
C7_246 n25_2 0 0.000092PF
C8_246 U280:A 0 0.000045PF
R1_246 U280:A n25_2 4.000000
R2_246 n25_2 n25_3 0.912000
R3_246 n25_3 n25_4 4.000000
R4_246 n25_5 n25_4 1.368000
R5_246 n25_5 n25_6 4.000000
R6_246 n25_6 n25_7 0.152000
R7_246 n25_7 clk_r_REG41_S2:Q 4.000000

C1_112 U264:Z 0 0.000045PF
C2_112 Q_PNN753_6 0 0.000121PF
C3_112 Q_PNN753_5 0 0.000141PF
C4_112 Q_PNN753_4 0 0.000141PF
C5_112 Q_PNN753_3 0 0.000136PF
C6_112 Q_PNN753_2 0 0.000136PF
C7_112 oDFF_30_q_reg:D 0 0.000045PF
R1_112 oDFF_30_q_reg:D Q_PNN753_2 4.000000
R2_112 Q_PNN753_2 Q_PNN753_3 1.368000
R3_112 Q_PNN753_3 Q_PNN753_4 4.000000
R4_112 Q_PNN753_5 Q_PNN753_4 1.216000
R5_112 Q_PNN753_5 Q_PNN753_6 4.000000
R6_112 Q_PNN753_6 U264:Z 4.000000

C1_290 U313:Z 0 0.000083PF
C2_290 n66_10 0 0.000106PF
C3_290 n66_9 0 0.000282PF
C4_290 n66_8 0 0.000282PF
C5_290 U203:B 0 0.000090PF
C6_290 n66_6 0 0.000135PF
C7_290 n66_5 0 0.000135PF
C8_290 n66_4 0 0.000292PF
C9_290 n66_3 0 0.000292PF
C10_290 n66_2 0 0.000121PF
C11_290 U201:B 0 0.000045PF
R1_290 U201:B n66_2 4.000000
R2_290 n66_2 n66_3 4.000000
R3_290 n66_4 n66_3 3.496000
R4_290 n66_4 n66_5 4.000000
R5_290 n66_6 n66_5 1.368000
R6_290 n66_6 U203:B 4.000000
R7_290 U203:B n66_8 4.000000
R8_290 n66_9 n66_8 3.496000
R9_290 n66_9 n66_10 4.000000
R10_290 U313:Z n66_10 0.760000

C1_148 U183:A 0 0.000045PF
C2_148 c0_n19_14 0 0.000054PF
C3_148 c0_n19_12 0 0.000125PF
C4_148 c0_n19_15 0 0.001174PF
C5_148 c0_n19_17 0 0.001174PF
C6_148 c0_n19_18 0 0.000112PF
C7_148 c0_n19_19 0 0.000112PF
C8_148 clk_r_REG27_S2:D 0 0.000045PF
C9_148 U256:Z 0 0.000045PF
C10_148 c0_n19_11 0 0.000039PF
C11_148 c0_n19_9 0 0.000055PF
C12_148 c0_n19_7 0 0.000741PF
C13_148 c0_n19_5 0 0.000741PF
C14_148 c0_n19_2 0 0.000072PF
C15_148 c0_n19_4 0 0.000057PF
C16_148 c0_n19_6 0 0.000181PF
C17_148 c0_n19_8 0 0.000181PF
C18_148 c0_n19_10 0 0.000089PF
C19_148 U181:A 0 0.000045PF
C20_148 c0_n19_1 0 0.000033PF
R1_148 c0_n19_2 c0_n19_1 0.152000
R2_148 c0_n19_1 U181:A 4.000000
R3_148 c0_n19_4 c0_n19_2 0.456000
R4_148 c0_n19_2 c0_n19_5 4.000000
R5_148 c0_n19_4 c0_n19_6 4.000000
R6_148 c0_n19_5 c0_n19_7 3.648000
R7_148 c0_n19_8 c0_n19_6 2.128000
R8_148 c0_n19_7 c0_n19_9 4.000000
R9_148 c0_n19_8 c0_n19_10 4.000000
R10_148 c0_n19_9 c0_n19_11 0.152000
R11_148 c0_n19_12 c0_n19_10 1.064000
R12_148 c0_n19_11 U256:Z 4.000000
R13_148 c0_n19_14 c0_n19_12 0.152000
R14_148 c0_n19_12 c0_n19_15 4.000000
R15_148 c0_n19_14 U183:A 4.000000
R16_148 c0_n19_17 c0_n19_15 3.800000
R17_148 c0_n19_17 c0_n19_18 4.000000
R18_148 c0_n19_18 c0_n19_19 1.824000
R19_148 c0_n19_19 clk_r_REG27_S2:D 4.000000

C1_211 U218:Z 0 0.000045PF
C2_211 n149_7 0 0.000135PF
C3_211 n149_6 0 0.000135PF
C4_211 n149_5 0 0.000697PF
C5_211 n149_4 0 0.000697PF
C6_211 n149_3 0 0.000100PF
C7_211 n149_2 0 0.000100PF
C8_211 U216:B 0 0.000045PF
R1_211 U216:B n149_2 4.000000
R2_211 n149_3 n149_2 0.760000
R3_211 n149_3 n149_4 4.000000
R4_211 n149_4 n149_5 1.976000
R5_211 n149_5 n149_6 4.000000
R6_211 n149_7 n149_6 1.368000
R7_211 n149_7 U218:Z 4.000000

C1_180 U258:Z 0 0.000045PF
C2_180 n115_7 0 0.000138PF
C3_180 n115_6 0 0.000138PF
C4_180 n115_5 0 0.000364PF
C5_180 n115_4 0 0.000364PF
C6_180 n115_3 0 0.000117PF
C7_180 n115_2 0 0.000117PF
C8_180 U256:B 0 0.000045PF
R1_180 U256:B n115_2 4.000000
R2_180 n115_3 n115_2 0.760000
R3_180 n115_3 n115_4 4.000000
R4_180 n115_4 n115_5 1.368000
R5_180 n115_5 n115_6 4.000000
R6_180 n115_7 n115_6 1.368000
R7_180 n115_7 U258:Z 4.000000

C1_205 U250:Z 0 0.000045PF
C2_205 n143_12 0 0.000121PF
C3_205 n143_11 0 0.000213PF
C4_205 n143_10 0 0.000213PF
C5_205 n143_9 0 0.000843PF
C6_205 n143_8 0 0.000843PF
C7_205 U220:A 0 0.000090PF
C8_205 n143_6 0 0.000047PF
C9_205 n143_5 0 0.000047PF
C10_205 n143_4 0 0.000487PF
C11_205 n143_3 0 0.000487PF
C12_205 n143_2 0 0.000121PF
C13_205 U208:B 0 0.000045PF
R1_205 U208:B n143_2 4.000000
R2_205 n143_2 n143_3 4.000000
R3_205 n143_3 n143_4 1.976000
R4_205 n143_4 n143_5 4.000000
R5_205 n143_6 n143_5 0.304000
R6_205 n143_6 U220:A 4.000000
R7_205 U220:A n143_8 4.000000
R8_205 n143_9 n143_8 7.600000
R9_205 n143_9 n143_10 4.000000
R10_205 n143_10 n143_11 1.976000
R11_205 n143_11 n143_12 4.000000
R12_205 n143_12 U250:Z 4.000000

C1_275 U312:A 0 0.000045PF
C2_275 n52_6 0 0.000121PF
C3_275 n52_5 0 0.000137PF
C4_275 n52_4 0 0.000137PF
C5_275 n52_3 0 0.000050PF
C6_275 n52_2 0 0.000034PF
C7_275 clk_r_REG13_S2:Q 0 0.000045PF
R1_275 clk_r_REG13_S2:Q n52_2 4.000000
R2_275 n52_2 n52_3 0.152000
R3_275 n52_3 n52_4 4.000000
R4_275 n52_4 n52_5 0.912000
R5_275 n52_5 n52_6 4.000000
R6_275 n52_6 U312:A 4.000000

C1_233 U264:A 0 0.000045PF
C2_233 n17_7 0 0.000045PF
C3_233 n17_6 0 0.000045PF
C4_233 n17_5 0 0.000296PF
C5_233 n17_4 0 0.000296PF
C6_233 n17_3 0 0.000137PF
C7_233 n17_2 0 0.000137PF
C8_233 clk_r_REG49_S2:Q 0 0.000045PF
R1_233 clk_r_REG49_S2:Q n17_2 4.000000
R2_233 n17_3 n17_2 1.672000
R3_233 n17_3 n17_4 4.000000
R4_233 n17_5 n17_4 1.216000
R5_233 n17_5 n17_6 4.000000
R6_233 n17_7 n17_6 0.456000
R7_233 n17_7 U264:A 4.000000

C1_174 U273:A 0 0.000045PF
C2_174 n11_5 0 0.000121PF
C3_174 n11_2 0 0.000270PF
C4_174 n11_4 0 0.000174PF
C5_174 n11_7 0 0.000121PF
C6_174 U265:A 0 0.000045PF
C7_174 clk_r_REG27_S2:Q 0 0.000045PF
C8_174 n11_6 0 0.000052PF
C9_174 n11_3 0 0.000052PF
C10_174 n11_1 0 0.000115PF
R1_174 n11_2 n11_1 1.976000
R2_174 n11_1 n11_3 4.000000
R3_174 n11_4 n11_2 1.672000
R4_174 n11_2 n11_5 4.000000
R5_174 n11_6 n11_3 0.304000
R6_174 n11_4 n11_7 4.000000
R7_174 n11_5 U273:A 4.000000
R8_174 n11_6 clk_r_REG27_S2:Q 4.000000
R9_174 n11_7 U265:A 4.000000

C1_78 PNN85 0 0.001985PF
C2_78 PNN85_5 0 0.002040PF
C3_78 PNN85_4 0 0.000580PF
C4_78 PNN85_3 0 0.000545PF
C5_78 PNN85_2 0 0.000121PF
C6_78 iDFF_22_q_reg:D 0 0.000045PF
R1_78 iDFF_22_q_reg:D PNN85_2 4.000000
R2_78 PNN85_2 PNN85_3 4.000000
R3_78 PNN85_3 PNN85_4 6.384000
R4_78 PNN85_5 PNN85_4 0.152000
R5_78 PNN85_5 PNN85 24.167999

C1_301 U264:B 0 0.000045PF
C2_301 n76_5 0 0.000121PF
C3_301 n76_4 0 0.000281PF
C4_301 n76_3 0 0.000281PF
C5_301 n76_2 0 0.000121PF
C6_301 U265:Z 0 0.000045PF
R1_301 U265:Z n76_2 4.000000
R2_301 n76_2 n76_3 4.000000
R3_301 n76_4 n76_3 1.976000
R4_301 n76_4 n76_5 4.000000
R5_301 n76_5 U264:B 4.000000

C1_181 U256:C 0 0.000045PF
C2_181 n116_7 0 0.000090PF
C3_181 n116_6 0 0.000090PF
C4_181 n116_5 0 0.000110PF
C5_181 n116_4 0 0.000110PF
C6_181 n116_3 0 0.000100PF
C7_181 n116_2 0 0.000100PF
C8_181 U257:Z 0 0.000045PF
R1_181 U257:Z n116_2 4.000000
R2_181 n116_3 n116_2 1.368000
R3_181 n116_3 n116_4 4.000000
R4_181 n116_4 n116_5 0.456000
R5_181 n116_5 n116_6 4.000000
R6_181 n116_7 n116_6 0.304000
R7_181 n116_7 U256:C 4.000000

C1_33 clk_r_REG37_S2:D 0 0.000045PF
C2_33 INP_PNN69_15 0 0.000041PF
C3_33 INP_PNN69_12 0 0.000041PF
C4_33 INP_PNN69_9 0 0.000207PF
C5_33 INP_PNN69_6 0 0.000481PF
C6_33 INP_PNN69_4 0 0.000322PF
C7_33 INP_PNN69_2 0 0.000418PF
C8_33 INP_PNN69_5 0 0.000428PF
C9_33 INP_PNN69_7 0 0.000428PF
C10_33 INP_PNN69_10 0 0.000052PF
C11_33 INP_PNN69_13 0 0.000035PF
C12_33 U259:B 0 0.000045PF
C13_33 iDFF_18_q_reg:Q 0 0.000045PF
C14_33 INP_PNN69_14 0 0.000055PF
C15_33 INP_PNN69_11 0 0.000071PF
C16_33 INP_PNN69_8 0 0.000292PF
C17_33 U254:B 0 0.000045PF
C18_33 INP_PNN69_1 0 0.000115PF
R1_33 INP_PNN69_2 INP_PNN69_1 1.216000
R2_33 INP_PNN69_1 U254:B 4.000000
R3_33 INP_PNN69_4 INP_PNN69_2 3.952000
R4_33 INP_PNN69_2 INP_PNN69_5 4.000000
R5_33 INP_PNN69_4 INP_PNN69_6 4.000000
R6_33 INP_PNN69_7 INP_PNN69_5 1.824000
R7_33 INP_PNN69_8 INP_PNN69_6 1.216000
R8_33 INP_PNN69_6 INP_PNN69_9 1.520000
R9_33 INP_PNN69_7 INP_PNN69_10 4.000000
R10_33 INP_PNN69_8 INP_PNN69_11 4.000000
R11_33 INP_PNN69_9 INP_PNN69_12 4.000000
R12_33 INP_PNN69_13 INP_PNN69_10 0.152000
R13_33 INP_PNN69_11 INP_PNN69_14 0.152000
R14_33 INP_PNN69_15 INP_PNN69_12 0.304000
R15_33 INP_PNN69_13 U259:B 4.000000
R16_33 INP_PNN69_14 iDFF_18_q_reg:Q 4.000000
R17_33 INP_PNN69_15 clk_r_REG37_S2:D 4.000000

C1_217 U208:Z 0 0.000045PF
C2_217 n155_7 0 0.000035PF
C3_217 n155_6 0 0.000051PF
C4_217 n155_5 0 0.000236PF
C5_217 n155_4 0 0.000236PF
C6_217 n155_3 0 0.000058PF
C7_217 n155_2 0 0.000041PF
C8_217 U160:B 0 0.000045PF
R1_217 U160:B n155_2 4.000000
R2_217 n155_3 n155_2 0.152000
R3_217 n155_3 n155_4 4.000000
R4_217 n155_4 n155_5 1.824000
R5_217 n155_5 n155_6 4.000000
R6_217 n155_7 n155_6 0.152000
R7_217 n155_7 U208:Z 4.000000

C1_147 U167:B 0 0.000045PF
C2_147 c0_n17_13 0 0.000060PF
C3_147 c0_n17_10 0 0.000060PF
C4_147 c0_n17_7 0 0.000757PF
C5_147 c0_n17_4 0 0.000665PF
C6_147 c0_n17_2 0 0.000186PF
C7_147 c0_n17_5 0 0.000129PF
C8_147 c0_n17_8 0 0.000129PF
C9_147 c0_n17_11 0 0.000371PF
C10_147 c0_n17_14 0 0.000371PF
C11_147 clk_r_REG15_S2:D 0 0.000045PF
C12_147 U177:A 0 0.000045PF
C13_147 c0_n17_15 0 0.000229PF
C14_147 c0_n17_12 0 0.000213PF
C15_147 c0_n17_9 0 0.000111PF
C16_147 U216:Z 0 0.000045PF
C17_147 c0_n17_21 0 0.000121PF
C18_147 c0_n17_20 0 0.000620PF
C19_147 c0_n17_18 0 0.000620PF
C20_147 U186:B 0 0.000045PF
C21_147 c0_n17_3 0 0.000086PF
C22_147 c0_n17_1 0 0.000220PF
R1_147 c0_n17_1 c0_n17_2 1.824000
R2_147 c0_n17_1 c0_n17_3 0.152000
R3_147 c0_n17_2 c0_n17_4 4.000000
R4_147 c0_n17_2 c0_n17_5 4.000000
R5_147 c0_n17_3 U186:B 4.000000
R6_147 c0_n17_4 c0_n17_7 2.888000
R7_147 c0_n17_8 c0_n17_5 1.064000
R8_147 c0_n17_7 c0_n17_9 1.520000
R9_147 c0_n17_7 c0_n17_10 4.000000
R10_147 c0_n17_8 c0_n17_11 4.000000
R11_147 c0_n17_9 c0_n17_12 4.000000
R12_147 c0_n17_10 c0_n17_13 0.304000
R13_147 c0_n17_11 c0_n17_14 2.280000
R14_147 c0_n17_15 c0_n17_12 1.824000
R15_147 c0_n17_13 U167:B 4.000000
R16_147 c0_n17_14 clk_r_REG15_S2:D 4.000000
R17_147 c0_n17_15 c0_n17_18 4.000000
R18_147 c0_n17_15 U177:A 4.000000
R19_147 c0_n17_18 c0_n17_20 1.824000
R20_147 c0_n17_20 c0_n17_21 4.000000
R21_147 c0_n17_21 U216:Z 4.000000

C1_182 U259:Z 0 0.000045PF
C2_182 n117_7 0 0.000306PF
C3_182 n117_6 0 0.000306PF
C4_182 n117_5 0 0.000902PF
C5_182 n117_4 0 0.000902PF
C6_182 n117_3 0 0.000046PF
C7_182 n117_2 0 0.000046PF
C8_182 U257:A 0 0.000045PF
R1_182 U257:A n117_2 4.000000
R2_182 n117_3 n117_2 0.304000
R3_182 n117_3 n117_4 4.000000
R4_182 n117_4 n117_5 6.840000
R5_182 n117_5 n117_6 4.000000
R6_182 n117_7 n117_6 1.368000
R7_182 n117_7 U259:Z 4.000000

C1_313 U283:Z 0 0.000045PF
C2_313 n87_5 0 0.000121PF
C3_313 n87_4 0 0.000108PF
C4_313 n87_3 0 0.000108PF
C5_313 n87_2 0 0.000121PF
C6_313 U282:B 0 0.000045PF
R1_313 U282:B n87_2 4.000000
R2_313 n87_2 n87_3 4.000000
R3_313 n87_4 n87_3 1.064000
R4_313 n87_4 n87_5 4.000000
R5_313 n87_5 U283:Z 4.000000

C1_237 U200:Z 0 0.000045PF
C2_237 n173_6 0 0.000588PF
C3_237 n173_5 0 0.000588PF
C4_237 n173_4 0 0.000232PF
C5_237 n173_3 0 0.000232PF
C6_237 n173_2 0 0.000121PF
C7_237 U199:A 0 0.000045PF
R1_237 U199:A n173_2 4.000000
R2_237 n173_2 n173_3 4.000000
R3_237 n173_4 n173_3 0.760000
R4_237 n173_4 n173_5 4.000000
R5_237 n173_5 n173_6 5.472000
R6_237 n173_6 U200:Z 4.000000

C1_289 U283:B 0 0.000045PF
C2_289 n65_11 0 0.000034PF
C3_289 n65_9 0 0.000050PF
C4_289 n65_7 0 0.000125PF
C5_289 n65_4 0 0.000125PF
C6_289 n65_2 0 0.000081PF
C7_289 U291:A 0 0.000045PF
C8_289 U312:Z 0 0.000045PF
C9_289 n65_10 0 0.000108PF
C10_289 n65_8 0 0.000108PF
C11_289 n65_6 0 0.000259PF
C12_289 n65_3 0 0.000259PF
C13_289 n65_1 0 0.000081PF
R1_289 n65_1 n65_2 0.760000
R2_289 n65_1 n65_3 4.000000
R3_289 n65_2 n65_4 4.000000
R4_289 n65_2 U291:A 4.000000
R5_289 n65_6 n65_3 2.432000
R6_289 n65_4 n65_7 1.976000
R7_289 n65_6 n65_8 4.000000
R8_289 n65_7 n65_9 4.000000
R9_289 n65_10 n65_8 1.216000
R10_289 n65_9 n65_11 0.152000
R11_289 n65_10 U312:Z 4.000000
R12_289 n65_11 U283:B 4.000000

C1_108 U272:Z 0 0.000045PF
C2_108 Q_PNN749_6 0 0.000121PF
C3_108 Q_PNN749_5 0 0.000674PF
C4_108 Q_PNN749_4 0 0.000674PF
C5_108 Q_PNN749_3 0 0.000127PF
C6_108 Q_PNN749_2 0 0.000127PF
C7_108 oDFF_26_q_reg:D 0 0.000045PF
R1_108 oDFF_26_q_reg:D Q_PNN749_2 4.000000
R2_108 Q_PNN749_3 Q_PNN749_2 1.520000
R3_108 Q_PNN749_3 Q_PNN749_4 4.000000
R4_108 Q_PNN749_4 Q_PNN749_5 3.800000
R5_108 Q_PNN749_5 Q_PNN749_6 4.000000
R6_108 Q_PNN749_6 U272:Z 4.000000

C1_242 U272:A 0 0.000045PF
C2_242 n21_5 0 0.000121PF
C3_242 n21_4 0 0.000117PF
C4_242 n21_3 0 0.000117PF
C5_242 n21_2 0 0.000121PF
C6_242 clk_r_REG45_S2:Q 0 0.000045PF
R1_242 clk_r_REG45_S2:Q n21_2 4.000000
R2_242 n21_2 n21_3 4.000000
R3_242 n21_4 n21_3 1.064000
R4_242 n21_4 n21_5 4.000000
R5_242 n21_5 U272:A 4.000000

C1_190 U171:B 0 0.000045PF
C2_190 n124_2 0 0.001493PF
C3_190 n124_4 0 0.000089PF
C4_190 n124_7 0 0.000139PF
C5_190 n124_9 0 0.000139PF
C6_190 n124_11 0 0.000055PF
C7_190 n124_13 0 0.000039PF
C8_190 U173:A 0 0.000090PF
C9_190 n124_15 0 0.000216PF
C10_190 n124_16 0 0.000216PF
C11_190 n124_17 0 0.000116PF
C12_190 n124_18 0 0.000116PF
C13_190 n124_19 0 0.000121PF
C14_190 U197:B 0 0.000045PF
C15_190 U214:Z 0 0.000045PF
C16_190 n124_10 0 0.000193PF
C17_190 n124_8 0 0.000193PF
C18_190 n124_6 0 0.000849PF
C19_190 n124_3 0 0.000849PF
C20_190 n124_1 0 0.001423PF
R1_190 n124_2 n124_1 12.768000
R2_190 n124_1 n124_3 4.000000
R3_190 n124_4 n124_2 1.064000
R4_190 n124_2 U171:B 4.000000
R5_190 n124_6 n124_3 3.496000
R6_190 n124_4 n124_7 4.000000
R7_190 n124_6 n124_8 4.000000
R8_190 n124_7 n124_9 0.456000
R9_190 n124_8 n124_10 1.368000
R10_190 n124_9 n124_11 4.000000
R11_190 n124_10 U214:Z 4.000000
R12_190 n124_13 n124_11 0.152000
R13_190 n124_13 U173:A 4.000000
R14_190 U173:A n124_15 4.000000
R15_190 n124_15 n124_16 1.976000
R16_190 n124_16 n124_17 4.000000
R17_190 n124_17 n124_18 1.368000
R18_190 n124_18 n124_19 4.000000
R19_190 n124_19 U197:B 4.000000

C1_103 U282:Z 0 0.000045PF
C2_103 Q_PNN744_6 0 0.000121PF
C3_103 Q_PNN744_5 0 0.000122PF
C4_103 Q_PNN744_4 0 0.000122PF
C5_103 Q_PNN744_3 0 0.000049PF
C6_103 Q_PNN744_2 0 0.000033PF
C7_103 oDFF_21_q_reg:D 0 0.000045PF
R1_103 oDFF_21_q_reg:D Q_PNN744_2 4.000000
R2_103 Q_PNN744_2 Q_PNN744_3 0.152000
R3_103 Q_PNN744_3 Q_PNN744_4 4.000000
R4_103 Q_PNN744_5 Q_PNN744_4 0.912000
R5_103 Q_PNN744_5 Q_PNN744_6 4.000000
R6_103 Q_PNN744_6 U282:Z 4.000000

C1_3 clk_r_REG45_S2:D 0 0.000045PF
C2_3 INP_PNN101_8 0 0.000310PF
C3_3 INP_PNN101_7 0 0.001542PF
C4_3 INP_PNN101_5 0 0.001542PF
C5_3 INP_PNN101_2 0 0.000246PF
C6_3 INP_PNN101_4 0 0.000218PF
C7_3 U214:C 0 0.000045PF
C8_3 iDFF_26_q_reg:Q 0 0.000045PF
C9_3 INP_PNN101_14 0 0.000035PF
C10_3 INP_PNN101_13 0 0.000051PF
C11_3 INP_PNN101_12 0 0.001216PF
C12_3 INP_PNN101_11 0 0.001216PF
C13_3 INP_PNN101_9 0 0.000310PF
C14_3 U257:C 0 0.000045PF
C15_3 INP_PNN101_1 0 0.000047PF
R1_3 INP_PNN101_1 INP_PNN101_2 0.304000
R2_3 INP_PNN101_1 U257:C 4.000000
R3_3 INP_PNN101_2 INP_PNN101_4 1.824000
R4_3 INP_PNN101_2 INP_PNN101_5 4.000000
R5_3 INP_PNN101_4 U214:C 4.000000
R6_3 INP_PNN101_7 INP_PNN101_5 9.272000
R7_3 INP_PNN101_7 INP_PNN101_8 4.000000
R8_3 INP_PNN101_8 INP_PNN101_9 1.216000
R9_3 INP_PNN101_8 clk_r_REG45_S2:D 4.000000
R10_3 INP_PNN101_9 INP_PNN101_11 4.000000
R11_3 INP_PNN101_12 INP_PNN101_11 4.712000
R12_3 INP_PNN101_12 INP_PNN101_13 4.000000
R13_3 INP_PNN101_13 INP_PNN101_14 0.152000
R14_3 INP_PNN101_14 iDFF_26_q_reg:Q 4.000000

C1_231 U160:Z 0 0.000045PF
C2_231 n168_7 0 0.000365PF
C3_231 n168_6 0 0.000365PF
C4_231 n168_5 0 0.000058PF
C5_231 n168_4 0 0.000058PF
C6_231 n168_3 0 0.000051PF
C7_231 n168_2 0 0.000051PF
C8_231 FE_OFCC1_n168:A 0 0.000045PF
R1_231 FE_OFCC1_n168:A n168_2 4.000000
R2_231 n168_3 n168_2 0.304000
R3_231 n168_3 n168_4 4.000000
R4_231 n168_4 n168_5 0.304000
R5_231 n168_5 n168_6 4.000000
R6_231 n168_7 n168_6 3.496000
R7_231 n168_7 U160:Z 4.000000

C1_208 U221:A 0 0.000045PF
C2_208 n146_7 0 0.000117PF
C3_208 n146_6 0 0.000117PF
C4_208 n146_5 0 0.000128PF
C5_208 n146_4 0 0.000128PF
C6_208 n146_3 0 0.000052PF
C7_208 n146_2 0 0.000036PF
C8_208 U223:Z 0 0.000045PF
R1_208 U223:Z n146_2 4.000000
R2_208 n146_3 n146_2 0.152000
R3_208 n146_3 n146_4 4.000000
R4_208 n146_5 n146_4 0.912000
R5_208 n146_5 n146_6 4.000000
R6_208 n146_7 n146_6 1.368000
R7_208 n146_7 U221:A 4.000000

C1_279 U166:B 0 0.000045PF
C2_279 n56_11 0 0.000337PF
C3_279 n56_10 0 0.000381PF
C4_279 n56_12 0 0.000641PF
C5_279 n56_15 0 0.000641PF
C6_279 n56_17 0 0.000121PF
C7_279 U164:B 0 0.000045PF
C8_279 U177:Z 0 0.000045PF
C9_279 n56_20 0 0.000121PF
C10_279 n56_18 0 0.000127PF
C11_279 n56_16 0 0.000127PF
C12_279 n56_13 0 0.000071PF
C13_279 U168:A 0 0.000045PF
C14_279 n56_5 0 0.000121PF
C15_279 n56_2 0 0.000443PF
C16_279 n56_4 0 0.000296PF
C17_279 n56_7 0 0.000099PF
C18_279 clk_r_REG16_S2:D 0 0.000045PF
C19_279 n56_6 0 0.000039PF
C20_279 n56_3 0 0.000055PF
C21_279 n56_1 0 0.000165PF
R1_279 n56_2 n56_1 0.760000
R2_279 n56_1 n56_3 4.000000
R3_279 n56_4 n56_2 1.064000
R4_279 n56_2 n56_5 4.000000
R5_279 n56_3 n56_6 0.152000
R6_279 n56_4 n56_7 4.000000
R7_279 n56_5 U168:A 4.000000
R8_279 n56_6 clk_r_REG16_S2:D 4.000000
R9_279 n56_10 n56_7 1.064000
R10_279 n56_11 n56_10 2.736000
R11_279 n56_10 n56_12 4.000000
R12_279 n56_13 n56_11 0.152000
R13_279 n56_11 U166:B 4.000000
R14_279 n56_15 n56_12 2.584000
R15_279 n56_13 n56_16 4.000000
R16_279 n56_15 n56_17 4.000000
R17_279 n56_16 n56_18 1.368000
R18_279 n56_17 U164:B 4.000000
R19_279 n56_18 n56_20 4.000000
R20_279 n56_20 U177:Z 4.000000

C1_32 U254:C 0 0.000045PF
C2_32 INP_PNN65_5 0 0.000147PF
C3_32 INP_PNN65_8 0 0.000695PF
C4_32 INP_PNN65_11 0 0.000695PF
C5_32 INP_PNN65_12 0 0.000121PF
C6_32 U221:B 0 0.000045PF
C7_32 iDFF_17_q_reg:Q 0 0.000045PF
C8_32 INP_PNN65_3 0 0.000130PF
C9_32 clk_r_REG36_S2:D 0 0.000045PF
C10_32 INP_PNN65_7 0 0.000046PF
C11_32 INP_PNN65_4 0 0.000046PF
C12_32 INP_PNN65_2 0 0.000099PF
C13_32 INP_PNN65_1 0 0.000099PF
R1_32 INP_PNN65_1 INP_PNN65_2 1.216000
R2_32 INP_PNN65_1 INP_PNN65_3 4.000000
R3_32 INP_PNN65_2 INP_PNN65_4 4.000000
R4_32 INP_PNN65_5 INP_PNN65_3 1.520000
R5_32 INP_PNN65_3 iDFF_17_q_reg:Q 4.000000
R6_32 INP_PNN65_4 INP_PNN65_7 0.304000
R7_32 INP_PNN65_5 INP_PNN65_8 4.000000
R8_32 INP_PNN65_5 U254:C 4.000000
R9_32 INP_PNN65_7 clk_r_REG36_S2:D 4.000000
R10_32 INP_PNN65_11 INP_PNN65_8 5.016000
R11_32 INP_PNN65_11 INP_PNN65_12 4.000000
R12_32 INP_PNN65_12 U221:B 4.000000

C1_251 clk_r_REG36_S2:Q 0 0.000045PF
C2_251 n30_6 0 0.000121PF
C3_251 n30_5 0 0.000129PF
C4_251 n30_4 0 0.000129PF
C5_251 n30_3 0 0.000049PF
C6_251 n30_2 0 0.000033PF
C7_251 U290:A 0 0.000045PF
R1_251 U290:A n30_2 4.000000
R2_251 n30_2 n30_3 0.152000
R3_251 n30_3 n30_4 4.000000
R4_251 n30_5 n30_4 1.368000
R5_251 n30_5 n30_6 4.000000
R6_251 n30_6 clk_r_REG36_S2:Q 4.000000

C1_319 U291:Z 0 0.000045PF
C2_319 n92_7 0 0.000120PF
C3_319 n92_6 0 0.000120PF
C4_319 n92_5 0 0.000092PF
C5_319 n92_4 0 0.000092PF
C6_319 n92_3 0 0.000071PF
C7_319 n92_2 0 0.000055PF
C8_319 U290:B 0 0.000045PF
R1_319 U290:B n92_2 4.000000
R2_319 n92_3 n92_2 0.152000
R3_319 n92_3 n92_4 4.000000
R4_319 n92_5 n92_4 0.608000
R5_319 n92_5 n92_6 4.000000
R6_319 n92_7 n92_6 1.368000
R7_319 n92_7 U291:Z 4.000000

C1_277 clk_r_REG16_S2:Q 0 0.000045PF
C2_277 n54_7 0 0.000260PF
C3_277 n54_6 0 0.000260PF
C4_277 n54_5 0 0.000437PF
C5_277 n54_4 0 0.000437PF
C6_277 n54_3 0 0.000076PF
C7_277 n54_2 0 0.000076PF
C8_277 U310:A 0 0.000045PF
R1_277 U310:A n54_2 4.000000
R2_277 n54_3 n54_2 0.456000
R3_277 n54_3 n54_4 4.000000
R4_277 n54_5 n54_4 3.496000
R5_277 n54_5 n54_6 4.000000
R6_277 n54_7 n54_6 1.064000
R7_277 n54_7 clk_r_REG16_S2:Q 4.000000

C1_36 iDFF_21_q_reg:Q 0 0.000045PF
C2_36 INP_PNN81_16 0 0.000033PF
C3_36 INP_PNN81_15 0 0.000049PF
C4_36 INP_PNN81_14 0 0.000622PF
C5_36 INP_PNN81_12 0 0.000622PF
C6_36 INP_PNN81_9 0 0.000197PF
C7_36 INP_PNN81_7 0 0.000132PF
C8_36 INP_PNN81_4 0 0.000512PF
C9_36 INP_PNN81_2 0 0.000586PF
C10_36 INP_PNN81_5 0 0.000171PF
C11_36 INP_PNN81_8 0 0.000171PF
C12_36 U212:C 0 0.000045PF
C13_36 clk_r_REG40_S2:D 0 0.000045PF
C14_36 INP_PNN81_11 0 0.000084PF
C15_36 U223:B 0 0.000045PF
C16_36 INP_PNN81_3 0 0.000121PF
C17_36 INP_PNN81_1 0 0.000092PF
R1_36 INP_PNN81_1 INP_PNN81_2 0.608000
R2_36 INP_PNN81_1 INP_PNN81_3 4.000000
R3_36 INP_PNN81_2 INP_PNN81_4 5.928000
R4_36 INP_PNN81_2 INP_PNN81_5 4.000000
R5_36 INP_PNN81_3 U223:B 4.000000
R6_36 INP_PNN81_4 INP_PNN81_7 4.000000
R7_36 INP_PNN81_8 INP_PNN81_5 1.976000
R8_36 INP_PNN81_7 INP_PNN81_9 1.368000
R9_36 INP_PNN81_8 U212:C 4.000000
R10_36 INP_PNN81_9 INP_PNN81_11 0.760000
R11_36 INP_PNN81_9 INP_PNN81_12 4.000000
R12_36 INP_PNN81_11 clk_r_REG40_S2:D 4.000000
R13_36 INP_PNN81_12 INP_PNN81_14 5.320000
R14_36 INP_PNN81_14 INP_PNN81_15 4.000000
R15_36 INP_PNN81_15 INP_PNN81_16 0.152000
R16_36 INP_PNN81_16 iDFF_21_q_reg:Q 4.000000

C1_238 U215:Z 0 0.000045PF
C2_238 n174_7 0 0.000280PF
C3_238 n174_6 0 0.000280PF
C4_238 n174_5 0 0.000178PF
C5_238 n174_4 0 0.000178PF
C6_238 n174_3 0 0.000368PF
C7_238 n174_2 0 0.000368PF
C8_238 U214:A 0 0.000045PF
R1_238 U214:A n174_2 4.000000
R2_238 n174_2 n174_3 1.520000
R3_238 n174_3 n174_4 4.000000
R4_238 n174_4 n174_5 0.608000
R5_238 n174_5 n174_6 4.000000
R6_238 n174_6 n174_7 1.976000
R7_238 n174_7 U215:Z 4.000000

C1_247 clk_r_REG40_S2:Q 0 0.000045PF
C2_247 n26_6 0 0.000121PF
C3_247 n26_5 0 0.000492PF
C4_247 n26_4 0 0.000492PF
C5_247 n26_3 0 0.000265PF
C6_247 n26_2 0 0.000265PF
C7_247 U282:A 0 0.000045PF
R1_247 U282:A n26_2 4.000000
R2_247 n26_2 n26_3 3.040000
R3_247 n26_3 n26_4 4.000000
R4_247 n26_5 n26_4 1.976000
R5_247 n26_5 n26_6 4.000000
R6_247 n26_6 clk_r_REG40_S2:Q 4.000000

C1_284 clk_r_REG24_S2:D 0 0.000045PF
C2_284 n60_16 0 0.000045PF
C3_284 n60_15 0 0.000045PF
C4_284 n60_14 0 0.000364PF
C5_284 n60_13 0 0.000364PF
C6_284 n60_12 0 0.000148PF
C7_284 n60_11 0 0.000148PF
C8_284 U182:Z 0 0.000090PF
C9_284 n60_8 0 0.000249PF
C10_284 n60_5 0 0.000249PF
C11_284 n60_2 0 0.000854PF
C12_284 n60_4 0 0.000685PF
C13_284 n60_7 0 0.000121PF
C14_284 U167:A 0 0.000045PF
C15_284 U164:A 0 0.000045PF
C16_284 n60_3 0 0.000121PF
C17_284 n60_1 0 0.000187PF
R1_284 n60_1 n60_2 0.608000
R2_284 n60_1 n60_3 4.000000
R3_284 n60_2 n60_4 1.824000
R4_284 n60_2 n60_5 4.000000
R5_284 n60_3 U164:A 4.000000
R6_284 n60_4 n60_7 4.000000
R7_284 n60_5 n60_8 1.216000
R8_284 n60_7 U167:A 4.000000
R9_284 n60_8 U182:Z 4.000000
R10_284 U182:Z n60_11 4.000000
R11_284 n60_11 n60_12 1.672000
R12_284 n60_12 n60_13 4.000000
R13_284 n60_14 n60_13 2.280000
R14_284 n60_14 n60_15 4.000000
R15_284 n60_15 n60_16 0.304000
R16_284 n60_16 clk_r_REG24_S2:D 4.000000

C1_99 oDFF_17_q_reg:D 0 0.000045PF
C2_99 Q_PNN740_7 0 0.000075PF
C3_99 Q_PNN740_6 0 0.000075PF
C4_99 Q_PNN740_5 0 0.000225PF
C5_99 Q_PNN740_4 0 0.000225PF
C6_99 Q_PNN740_3 0 0.000153PF
C7_99 Q_PNN740_2 0 0.000153PF
C8_99 U290:Z 0 0.000045PF
R1_99 U290:Z Q_PNN740_2 4.000000
R2_99 Q_PNN740_2 Q_PNN740_3 1.520000
R3_99 Q_PNN740_3 Q_PNN740_4 4.000000
R4_99 Q_PNN740_4 Q_PNN740_5 0.912000
R5_99 Q_PNN740_5 Q_PNN740_6 4.000000
R6_99 Q_PNN740_6 Q_PNN740_7 0.456000
R7_99 Q_PNN740_7 oDFF_17_q_reg:D 4.000000

C1_302 U267:Z 0 0.000045PF
C2_302 n77_5 0 0.000121PF
C3_302 n77_4 0 0.000445PF
C4_302 n77_3 0 0.000445PF
C5_302 n77_2 0 0.000121PF
C6_302 U266:B 0 0.000045PF
R1_302 U266:B n77_2 4.000000
R2_302 n77_2 n77_3 4.000000
R3_302 n77_3 n77_4 3.344000
R4_302 n77_4 n77_5 4.000000
R5_302 n77_5 U267:Z 4.000000

C1_306 U271:Z 0 0.000045PF
C2_306 n80_5 0 0.000121PF
C3_306 n80_4 0 0.000834PF
C4_306 n80_3 0 0.000834PF
C5_306 n80_2 0 0.000121PF
C6_306 U270:B 0 0.000045PF
R1_306 U270:B n80_2 4.000000
R2_306 n80_2 n80_3 4.000000
R3_306 n80_4 n80_3 4.864000
R4_306 n80_4 n80_5 4.000000
R5_306 n80_5 U271:Z 4.000000

C1_214 U219:Z 0 0.000045PF
C2_214 n151_5 0 0.000121PF
C3_214 n151_4 0 0.001856PF
C4_214 n151_3 0 0.001856PF
C5_214 n151_2 0 0.000121PF
C6_214 U217:A 0 0.000045PF
R1_214 U217:A n151_2 4.000000
R2_214 n151_2 n151_3 4.000000
R3_214 n151_3 n151_4 8.056000
R4_214 n151_4 n151_5 4.000000
R5_214 n151_5 U219:Z 4.000000

C1_195 U275:A 0 0.000045PF
C2_195 n13_9 0 0.000120PF
C3_195 n13_8 0 0.000120PF
C4_195 U267:A 0 0.000090PF
C5_195 n13_6 0 0.000121PF
C6_195 n13_5 0 0.000125PF
C7_195 n13_4 0 0.000125PF
C8_195 n13_3 0 0.000397PF
C9_195 n13_2 0 0.000397PF
C10_195 clk_r_REG12_S2:Q 0 0.000045PF
R1_195 clk_r_REG12_S2:Q n13_2 4.000000
R2_195 n13_2 n13_3 1.672000
R3_195 n13_3 n13_4 4.000000
R4_195 n13_5 n13_4 0.912000
R5_195 n13_5 n13_6 4.000000
R6_195 n13_6 U267:A 4.000000
R7_195 U267:A n13_8 4.000000
R8_195 n13_8 n13_9 1.216000
R9_195 n13_9 U275:A 4.000000

C1_185 clk_r_REG15_S2:Q 0 0.000045PF
C2_185 n12_9 0 0.000104PF
C3_185 n12_8 0 0.000104PF
C4_185 n12_7 0 0.000395PF
C5_185 n12_6 0 0.000395PF
C6_185 n12_5 0 0.000121PF
C7_185 U271:A 0 0.000090PF
C8_185 n12_3 0 0.000122PF
C9_185 n12_2 0 0.000122PF
C10_185 U263:A 0 0.000045PF
R1_185 U263:A n12_2 4.000000
R2_185 n12_3 n12_2 1.216000
R3_185 n12_3 U271:A 4.000000
R4_185 U271:A n12_5 4.000000
R5_185 n12_5 n12_6 4.000000
R6_185 n12_6 n12_7 1.672000
R7_185 n12_7 n12_8 4.000000
R8_185 n12_9 n12_8 1.672000
R9_185 n12_9 clk_r_REG15_S2:Q 4.000000

C1_77 PNN81 0 0.003498PF
C2_77 PNN81_3 0 0.003519PF
C3_77 PNN81_2 0 0.000121PF
C4_77 iDFF_21_q_reg:D 0 0.000045PF
R1_77 iDFF_21_q_reg:D PNN81_2 4.000000
R2_77 PNN81_2 PNN81_3 4.000000
R3_77 PNN81_3 PNN81 30.551999

C1_239 clk_r_REG48_S2:Q 0 0.000045PF
C2_239 n18_6 0 0.000121PF
C3_239 n18_5 0 0.000107PF
C4_239 n18_4 0 0.000107PF
C5_239 n18_3 0 0.000055PF
C6_239 n18_2 0 0.000039PF
C7_239 U266:A 0 0.000045PF
R1_239 U266:A n18_2 4.000000
R2_239 n18_3 n18_2 0.152000
R3_239 n18_3 n18_4 4.000000
R4_239 n18_4 n18_5 0.912000
R5_239 n18_5 n18_6 4.000000
R6_239 n18_6 clk_r_REG48_S2:Q 4.000000

C1_4 U217:C 0 0.000045PF
C2_4 INP_PNN105_10 0 0.000216PF
C3_4 INP_PNN105_11 0 0.000146PF
C4_4 INP_PNN105_13 0 0.000163PF
C5_4 INP_PNN105_14 0 0.000128PF
C6_4 U214:B 0 0.000045PF
C7_4 iDFF_27_q_reg:Q 0 0.000045PF
C8_4 INP_PNN105_5 0 0.000121PF
C9_4 INP_PNN105_2 0 0.000953PF
C10_4 INP_PNN105_4 0 0.000322PF
C11_4 INP_PNN105_7 0 0.000123PF
C12_4 clk_r_REG46_S2:D 0 0.000045PF
C13_4 INP_PNN105_6 0 0.000034PF
C14_4 INP_PNN105_3 0 0.000050PF
C15_4 INP_PNN105_1 0 0.000650PF
R1_4 INP_PNN105_1 INP_PNN105_2 2.584000
R2_4 INP_PNN105_1 INP_PNN105_3 4.000000
R3_4 INP_PNN105_2 INP_PNN105_4 1.368000
R4_4 INP_PNN105_2 INP_PNN105_5 4.000000
R5_4 INP_PNN105_6 INP_PNN105_3 0.152000
R6_4 INP_PNN105_4 INP_PNN105_7 4.000000
R7_4 INP_PNN105_5 iDFF_27_q_reg:Q 4.000000
R8_4 INP_PNN105_6 clk_r_REG46_S2:D 4.000000
R9_4 INP_PNN105_10 INP_PNN105_7 0.456000
R10_4 INP_PNN105_11 INP_PNN105_10 0.912000
R11_4 INP_PNN105_10 U217:C 4.000000
R12_4 INP_PNN105_13 INP_PNN105_11 0.152000
R13_4 INP_PNN105_14 INP_PNN105_13 0.912000
R14_4 INP_PNN105_14 U214:B 4.000000

C1_287 U310:Z 0 0.000045PF
C2_287 n63_2 0 0.000178PF
C3_287 n63_4 0 0.000289PF
C4_287 n63_6 0 0.000289PF
C5_287 n63_7 0 0.000121PF
C6_287 U287:A 0 0.000045PF
C7_287 U279:B 0 0.000045PF
C8_287 n63_1 0 0.000178PF
R1_287 n63_2 n63_1 1.064000
R2_287 n63_1 U279:B 4.000000
R3_287 n63_2 n63_4 4.000000
R4_287 n63_2 U310:Z 4.000000
R5_287 n63_4 n63_6 2.280000
R6_287 n63_6 n63_7 4.000000
R7_287 n63_7 U287:A 4.000000

C1_276 U309:A 0 0.000045PF
C2_276 n53_6 0 0.000121PF
C3_276 n53_5 0 0.000121PF
C4_276 n53_4 0 0.000111PF
C5_276 n53_3 0 0.000111PF
C6_276 n53_2 0 0.000121PF
C7_276 clk_r_REG25_S2:Q 0 0.000045PF
R1_276 clk_r_REG25_S2:Q n53_2 4.000000
R2_276 n53_2 n53_3 4.000000
R3_276 n53_4 n53_3 0.760000
R4_276 n53_4 n53_5 4.000000
R5_276 n53_5 n53_6 1.368000
R6_276 n53_6 U309:A 4.000000

C1_131 oDFF_17_q_reg:Q 0 0.000045PF
C2_131 Qout_PNN740_4 0 0.000033PF
C3_131 Qout_PNN740_3 0 0.000049PF
C4_131 Qout_PNN740_2 0 0.003824PF
C5_131 Qout_PNN740 0 0.003803PF
R1_131 Qout_PNN740_2 Qout_PNN740 33.287999
R2_131 Qout_PNN740_2 Qout_PNN740_3 4.000000
R3_131 Qout_PNN740_4 Qout_PNN740_3 0.152000
R4_131 Qout_PNN740_4 oDFF_17_q_reg:Q 4.000000

C1_109 oDFF_27_q_reg:D 0 0.000045PF
C2_109 Q_PNN750_7 0 0.000118PF
C3_109 Q_PNN750_6 0 0.000118PF
C4_109 Q_PNN750_5 0 0.000193PF
C5_109 Q_PNN750_4 0 0.000193PF
C6_109 Q_PNN750_3 0 0.000045PF
C7_109 Q_PNN750_2 0 0.000045PF
C8_109 U270:Z 0 0.000045PF
R1_109 U270:Z Q_PNN750_2 4.000000
R2_109 Q_PNN750_2 Q_PNN750_3 0.304000
R3_109 Q_PNN750_3 Q_PNN750_4 4.000000
R4_109 Q_PNN750_4 Q_PNN750_5 0.912000
R5_109 Q_PNN750_5 Q_PNN750_6 4.000000
R6_109 Q_PNN750_6 Q_PNN750_7 1.216000
R7_109 Q_PNN750_7 oDFF_27_q_reg:D 4.000000

C1_305 U261:A 0 0.000045PF
C2_305 n8_2 0 0.000050PF
C3_305 n8_4 0 0.000182PF
C4_305 n8_7 0 0.000182PF
C5_305 n8_9 0 0.000121PF
C6_305 U269:A 0 0.000045PF
C7_305 clk_r_REG24_S2:Q 0 0.000045PF
C8_305 n8_6 0 0.000058PF
C9_305 n8_3 0 0.000093PF
C10_305 n8_1 0 0.000085PF
R1_305 n8_1 n8_2 0.608000
R2_305 n8_3 n8_1 0.152000
R3_305 n8_2 n8_4 4.000000
R4_305 n8_2 U261:A 4.000000
R5_305 n8_6 n8_3 0.608000
R6_305 n8_4 n8_7 1.368000
R7_305 n8_6 clk_r_REG24_S2:Q 4.000000
R8_305 n8_7 n8_9 4.000000
R9_305 n8_9 U269:A 4.000000

C1_249 clk_r_REG38_S2:Q 0 0.000045PF
C2_249 n28_5 0 0.000121PF
C3_249 n28_4 0 0.000563PF
C4_249 n28_3 0 0.000563PF
C5_249 n28_2 0 0.000121PF
C6_249 U286:A 0 0.000045PF
R1_249 U286:A n28_2 4.000000
R2_249 n28_2 n28_3 4.000000
R3_249 n28_3 n28_4 2.432000
R4_249 n28_4 n28_5 4.000000
R5_249 n28_5 clk_r_REG38_S2:Q 4.000000

C1_310 U277:A 0 0.000045PF
C2_310 n84_13 0 0.000375PF
C3_310 n84_11 0 0.000711PF
C4_310 n84_9 0 0.000745PF
C5_310 n84_7 0 0.000905PF
C6_310 n84_4 0 0.000870PF
C7_310 n84_2 0 0.000247PF
C8_310 U279:A 0 0.000045PF
C9_310 U283:A 0 0.000078PF
C10_310 n84_15 0 0.000375PF
C11_310 U281:A 0 0.000045PF
C12_310 n84_24 0 0.000289PF
C13_310 n84_22 0 0.000289PF
C14_310 n84_20 0 0.000068PF
C15_310 U201:Z 0 0.000045PF
C16_310 n84_21 0 0.000513PF
C17_310 n84_19 0 0.000513PF
C18_310 n84_17 0 0.000130PF
C19_310 n84_14 0 0.000165PF
C20_310 n84_12 0 0.001836PF
C21_310 n84_10 0 0.001801PF
C22_310 n84_8 0 0.000121PF
C23_310 n84_6 0 0.000134PF
C24_310 n84_3 0 0.000134PF
C25_310 n84_1 0 0.000184PF
R1_310 n84_1 n84_2 1.216000
R2_310 n84_1 n84_3 4.000000
R3_310 n84_2 n84_4 4.000000
R4_310 n84_2 U279:A 4.000000
R5_310 n84_6 n84_3 0.912000
R6_310 n84_4 n84_7 6.080000
R7_310 n84_6 n84_8 4.000000
R8_310 n84_9 n84_7 0.152000
R9_310 n84_8 n84_10 4.000000
R10_310 n84_9 n84_11 8.664000
R11_310 n84_12 n84_10 12.616000
R12_310 n84_11 n84_13 4.000000
R13_310 n84_14 n84_12 0.152000
R14_310 n84_15 n84_13 5.168000
R15_310 n84_13 U277:A 4.000000
R16_310 n84_17 n84_14 0.912000
R17_310 n84_15 U283:A 4.000000
R18_310 n84_17 n84_19 4.000000
R19_310 U283:A n84_20 0.456000
R20_310 n84_21 n84_19 5.928000
R21_310 n84_20 n84_22 4.000000
R22_310 n84_21 U201:Z 4.000000
R23_310 n84_24 n84_22 3.952000
R24_310 n84_24 U281:A 4.000000

C1_41 clk_r_REG44_S2:D 0 0.000045PF
C2_41 INP_PNN97_10 0 0.000121PF
C3_41 INP_PNN97_8 0 0.000289PF
C4_41 INP_PNN97_6 0 0.000289PF
C5_41 INP_PNN97_4 0 0.000121PF
C6_41 U223:A 0 0.000199PF
C7_41 iDFF_25_q_reg:Q 0 0.000244PF
C8_41 INP_PNN97_11 0 0.000218PF
C9_41 INP_PNN97_9 0 0.000218PF
C10_41 INP_PNN97_7 0 0.001050PF
C11_41 INP_PNN97_5 0 0.001050PF
C12_41 INP_PNN97_3 0 0.000245PF
C13_41 INP_PNN97_2 0 0.000245PF
C14_41 U215:A 0 0.000090PF
R1_41 U215:A INP_PNN97_2 4.000000
R2_41 INP_PNN97_3 INP_PNN97_2 2.432000
R3_41 U215:A INP_PNN97_4 4.000000
R4_41 INP_PNN97_3 INP_PNN97_5 4.000000
R5_41 INP_PNN97_4 INP_PNN97_6 4.000000
R6_41 INP_PNN97_5 INP_PNN97_7 4.408000
R7_41 INP_PNN97_8 INP_PNN97_6 3.800000
R8_41 INP_PNN97_7 INP_PNN97_9 4.000000
R9_41 INP_PNN97_8 INP_PNN97_10 4.000000
R10_41 INP_PNN97_11 INP_PNN97_9 1.672000
R11_41 INP_PNN97_10 clk_r_REG44_S2:D 4.000000
R12_41 INP_PNN97_11 iDFF_25_q_reg:Q 4.000000
R13_41 iDFF_25_q_reg:Q U223:A 1.976000

C1_34 clk_r_REG38_S2:D 0 0.000069PF
C2_34 INP_PNN73_17 0 0.000091PF
C3_34 INP_PNN73_16 0 0.000121PF
C4_34 INP_PNN73_15 0 0.000092PF
C5_34 INP_PNN73_14 0 0.000092PF
C6_34 INP_PNN73_13 0 0.000071PF
C7_34 INP_PNN73_12 0 0.000055PF
C8_34 U255:B 0 0.000090PF
C9_34 INP_PNN73_10 0 0.000240PF
C10_34 INP_PNN73_9 0 0.000240PF
C11_34 iDFF_19_q_reg:Q 0 0.000090PF
C12_34 INP_PNN73_7 0 0.000034PF
C13_34 INP_PNN73_6 0 0.000050PF
C14_34 INP_PNN73_5 0 0.000292PF
C15_34 INP_PNN73_4 0 0.000292PF
C16_34 INP_PNN73_3 0 0.000049PF
C17_34 INP_PNN73_2 0 0.000033PF
C18_34 U219:B 0 0.000045PF
R1_34 U219:B INP_PNN73_2 4.000000
R2_34 INP_PNN73_3 INP_PNN73_2 0.152000
R3_34 INP_PNN73_3 INP_PNN73_4 4.000000
R4_34 INP_PNN73_4 INP_PNN73_5 3.192000
R5_34 INP_PNN73_5 INP_PNN73_6 4.000000
R6_34 INP_PNN73_7 INP_PNN73_6 0.152000
R7_34 INP_PNN73_7 iDFF_19_q_reg:Q 4.000000
R8_34 iDFF_19_q_reg:Q INP_PNN73_9 4.000000
R9_34 INP_PNN73_9 INP_PNN73_10 1.672000
R10_34 INP_PNN73_10 U255:B 4.000000
R11_34 U255:B INP_PNN73_12 4.000000
R12_34 INP_PNN73_13 INP_PNN73_12 0.152000
R13_34 INP_PNN73_13 INP_PNN73_14 4.000000
R14_34 INP_PNN73_15 INP_PNN73_14 0.760000
R15_34 INP_PNN73_15 INP_PNN73_16 4.000000
R16_34 INP_PNN73_16 INP_PNN73_17 4.000000
R17_34 clk_r_REG38_S2:D INP_PNN73_17 0.760000

C1_288 U309:Z 0 0.000045PF
C2_288 n64_6 0 0.000121PF
C3_288 n64_5 0 0.000343PF
C4_288 n64_4 0 0.000343PF
C5_288 n64_3 0 0.000121PF
C6_288 U285:A 0 0.000183PF
C7_288 U277:B 0 0.000138PF
R1_288 U285:A U277:B 1.368000
R2_288 U285:A n64_3 4.000000
R3_288 n64_3 n64_4 4.000000
R4_288 n64_5 n64_4 2.736000
R5_288 n64_5 n64_6 4.000000
R6_288 n64_6 U309:Z 4.000000

C1_106 U276:Z 0 0.000045PF
C2_106 Q_PNN747_5 0 0.000121PF
C3_106 Q_PNN747_4 0 0.000238PF
C4_106 Q_PNN747_3 0 0.000238PF
C5_106 Q_PNN747_2 0 0.000121PF
C6_106 oDFF_24_q_reg:D 0 0.000045PF
R1_106 oDFF_24_q_reg:D Q_PNN747_2 4.000000
R2_106 Q_PNN747_2 Q_PNN747_3 4.000000
R3_106 Q_PNN747_4 Q_PNN747_3 0.912000
R4_106 Q_PNN747_4 Q_PNN747_5 4.000000
R5_106 Q_PNN747_5 U276:Z 4.000000

C1_303 U269:Z 0 0.000045PF
C2_303 n78_6 0 0.000121PF
C3_303 n78_5 0 0.000396PF
C4_303 n78_4 0 0.000396PF
C5_303 n78_3 0 0.000171PF
C6_303 n78_2 0 0.000171PF
C7_303 U268:B 0 0.000045PF
R1_303 U268:B n78_2 4.000000
R2_303 n78_3 n78_2 1.824000
R3_303 n78_3 n78_4 4.000000
R4_303 n78_5 n78_4 4.408000
R5_303 n78_5 n78_6 4.000000
R6_303 n78_6 U269:Z 4.000000

C1_309 U277:Z 0 0.000045PF
C2_309 n83_5 0 0.000121PF
C3_309 n83_4 0 0.000108PF
C4_309 n83_3 0 0.000108PF
C5_309 n83_2 0 0.000121PF
C6_309 U276:B 0 0.000045PF
R1_309 U276:B n83_2 4.000000
R2_309 n83_2 n83_3 4.000000
R3_309 n83_4 n83_3 1.064000
R4_309 n83_4 n83_5 4.000000
R5_309 n83_5 U277:Z 4.000000

C1_244 clk_r_REG43_S2:Q 0 0.000045PF
C2_244 n23_7 0 0.000136PF
C3_244 n23_6 0 0.000136PF
C4_244 n23_5 0 0.000284PF
C5_244 n23_4 0 0.000284PF
C6_244 n23_3 0 0.000039PF
C7_244 n23_2 0 0.000039PF
C8_244 U276:A 0 0.000045PF
R1_244 U276:A n23_2 4.000000
R2_244 n23_2 n23_3 0.304000
R3_244 n23_3 n23_4 4.000000
R4_244 n23_4 n23_5 2.280000
R5_244 n23_5 n23_6 4.000000
R6_244 n23_6 n23_7 1.520000
R7_244 n23_7 clk_r_REG43_S2:Q 4.000000

C1_101 U286:Z 0 0.000045PF
C2_101 Q_PNN742_7 0 0.000033PF
C3_101 Q_PNN742_6 0 0.000050PF
C4_101 Q_PNN742_5 0 0.000159PF
C5_101 Q_PNN742_4 0 0.000159PF
C6_101 Q_PNN742_3 0 0.000147PF
C7_101 Q_PNN742_2 0 0.000147PF
C8_101 oDFF_19_q_reg:D 0 0.000045PF
R1_101 oDFF_19_q_reg:D Q_PNN742_2 4.000000
R2_101 Q_PNN742_3 Q_PNN742_2 1.824000
R3_101 Q_PNN742_3 Q_PNN742_4 4.000000
R4_101 Q_PNN742_5 Q_PNN742_4 1.520000
R5_101 Q_PNN742_5 Q_PNN742_6 4.000000
R6_101 Q_PNN742_7 Q_PNN742_6 0.152000
R7_101 Q_PNN742_7 U286:Z 4.000000

C1_243 clk_r_REG44_S2:Q 0 0.000045PF
C2_243 n22_7 0 0.000135PF
C3_243 n22_6 0 0.000135PF
C4_243 n22_5 0 0.000685PF
C5_243 n22_4 0 0.000685PF
C6_243 n22_3 0 0.000081PF
C7_243 n22_2 0 0.000081PF
C8_243 U274:A 0 0.000045PF
R1_243 U274:A n22_2 4.000000
R2_243 n22_3 n22_2 0.760000
R3_243 n22_3 n22_4 4.000000
R4_243 n22_4 n22_5 8.360000
R5_243 n22_5 n22_6 4.000000
R6_243 n22_7 n22_6 1.368000
R7_243 n22_7 clk_r_REG44_S2:Q 4.000000

C1_35 clk_r_REG39_S2:D 0 0.000045PF
C2_35 INP_PNN77_9 0 0.000082PF
C3_35 INP_PNN77_8 0 0.000045PF
C4_35 INP_PNN77_7 0 0.000200PF
C5_35 INP_PNN77_5 0 0.000200PF
C6_35 INP_PNN77_2 0 0.000323PF
C7_35 INP_PNN77_4 0 0.000308PF
C8_35 U255:A 0 0.000045PF
C9_35 iDFF_20_q_reg:Q 0 0.000045PF
C10_35 INP_PNN77_13 0 0.000069PF
C11_35 INP_PNN77_12 0 0.000104PF
C12_35 INP_PNN77_10 0 0.000090PF
C13_35 U209:B 0 0.000045PF
C14_35 INP_PNN77_1 0 0.000033PF
R1_35 INP_PNN77_2 INP_PNN77_1 0.152000
R2_35 INP_PNN77_1 U209:B 4.000000
R3_35 INP_PNN77_4 INP_PNN77_2 2.280000
R4_35 INP_PNN77_2 INP_PNN77_5 4.000000
R5_35 INP_PNN77_4 U255:A 4.000000
R6_35 INP_PNN77_5 INP_PNN77_7 1.520000
R7_35 INP_PNN77_7 INP_PNN77_8 4.000000
R8_35 INP_PNN77_8 INP_PNN77_9 0.456000
R9_35 INP_PNN77_9 INP_PNN77_10 0.760000
R10_35 INP_PNN77_9 clk_r_REG39_S2:D 4.000000
R11_35 INP_PNN77_10 INP_PNN77_12 0.152000
R12_35 INP_PNN77_12 INP_PNN77_13 0.608000
R13_35 INP_PNN77_13 iDFF_20_q_reg:Q 4.000000

C1_300 U263:Z 0 0.000045PF
C2_300 n75_6 0 0.000171PF
C3_300 n75_5 0 0.000171PF
C4_300 n75_4 0 0.000123PF
C5_300 n75_3 0 0.000123PF
C6_300 n75_2 0 0.000121PF
C7_300 U262:B 0 0.000045PF
R1_300 U262:B n75_2 4.000000
R2_300 n75_2 n75_3 4.000000
R3_300 n75_4 n75_3 0.456000
R4_300 n75_4 n75_5 4.000000
R5_300 n75_6 n75_5 1.824000
R6_300 n75_6 U263:Z 4.000000

C1_113 U262:Z 0 0.000045PF
C2_113 Q_PNN754_6 0 0.000121PF
C3_113 Q_PNN754_5 0 0.000070PF
C4_113 Q_PNN754_4 0 0.000070PF
C5_113 Q_PNN754_3 0 0.000142PF
C6_113 Q_PNN754_2 0 0.000142PF
C7_113 oDFF_31_q_reg:D 0 0.000045PF
R1_113 oDFF_31_q_reg:D Q_PNN754_2 4.000000
R2_113 Q_PNN754_3 Q_PNN754_2 1.520000
R3_113 Q_PNN754_3 Q_PNN754_4 4.000000
R4_113 Q_PNN754_5 Q_PNN754_4 0.608000
R5_113 Q_PNN754_5 Q_PNN754_6 4.000000
R6_113 Q_PNN754_6 U262:Z 4.000000

C1_240 U268:A 0 0.000045PF
C2_240 n19_5 0 0.000121PF
C3_240 n19_4 0 0.000079PF
C4_240 n19_3 0 0.000079PF
C5_240 n19_2 0 0.000121PF
C6_240 clk_r_REG47_S2:Q 0 0.000045PF
R1_240 clk_r_REG47_S2:Q n19_2 4.000000
R2_240 n19_2 n19_3 4.000000
R3_240 n19_4 n19_3 0.760000
R4_240 n19_4 n19_5 4.000000
R5_240 n19_5 U268:A 4.000000

C1_5 U207:C 0 0.000045PF
C2_5 INP_PNN109_17 0 0.000038PF
C3_5 INP_PNN109_16 0 0.000055PF
C4_5 INP_PNN109_15 0 0.000201PF
C5_5 INP_PNN109_14 0 0.000201PF
C6_5 INP_PNN109_13 0 0.000050PF
C7_5 INP_PNN109_12 0 0.000034PF
C8_5 iDFF_28_q_reg:Q 0 0.000090PF
C9_5 INP_PNN109_7 0 0.000121PF
C10_5 INP_PNN109_4 0 0.000132PF
C11_5 INP_PNN109_2 0 0.000320PF
C12_5 INP_PNN109_5 0 0.000162PF
C13_5 INP_PNN109_8 0 0.000162PF
C14_5 U215:B 0 0.000045PF
C15_5 clk_r_REG47_S2:D 0 0.000045PF
C16_5 INP_PNN109_6 0 0.000035PF
C17_5 INP_PNN109_3 0 0.000052PF
C18_5 INP_PNN109_1 0 0.000206PF
R1_5 INP_PNN109_1 INP_PNN109_2 1.520000
R2_5 INP_PNN109_1 INP_PNN109_3 4.000000
R3_5 INP_PNN109_2 INP_PNN109_4 0.912000
R4_5 INP_PNN109_2 INP_PNN109_5 4.000000
R5_5 INP_PNN109_6 INP_PNN109_3 0.152000
R6_5 INP_PNN109_4 INP_PNN109_7 4.000000
R7_5 INP_PNN109_8 INP_PNN109_5 2.432000
R8_5 INP_PNN109_6 clk_r_REG47_S2:D 4.000000
R9_5 INP_PNN109_7 iDFF_28_q_reg:Q 4.000000
R10_5 INP_PNN109_8 U215:B 4.000000
R11_5 iDFF_28_q_reg:Q INP_PNN109_12 4.000000
R12_5 INP_PNN109_12 INP_PNN109_13 0.152000
R13_5 INP_PNN109_13 INP_PNN109_14 4.000000
R14_5 INP_PNN109_14 INP_PNN109_15 1.216000
R15_5 INP_PNN109_15 INP_PNN109_16 4.000000
R16_5 INP_PNN109_16 INP_PNN109_17 0.152000
R17_5 INP_PNN109_17 U207:C 4.000000

C1_248 clk_r_REG39_S2:Q 0 0.000045PF
C2_248 n27_6 0 0.000121PF
C3_248 n27_5 0 0.000375PF
C4_248 n27_4 0 0.000375PF
C5_248 n27_3 0 0.000055PF
C6_248 n27_2 0 0.000039PF
C7_248 U284:A 0 0.000045PF
R1_248 U284:A n27_2 4.000000
R2_248 n27_3 n27_2 0.152000
R3_248 n27_3 n27_4 4.000000
R4_248 n27_5 n27_4 1.368000
R5_248 n27_5 n27_6 4.000000
R6_248 n27_6 clk_r_REG39_S2:Q 4.000000

C1_110 U268:Z 0 0.000045PF
C2_110 Q_PNN751_7 0 0.000047PF
C3_110 Q_PNN751_6 0 0.000047PF
C4_110 Q_PNN751_5 0 0.000110PF
C5_110 Q_PNN751_4 0 0.000110PF
C6_110 Q_PNN751_3 0 0.000152PF
C7_110 Q_PNN751_2 0 0.000152PF
C8_110 oDFF_28_q_reg:D 0 0.000045PF
R1_110 oDFF_28_q_reg:D Q_PNN751_2 4.000000
R2_110 Q_PNN751_3 Q_PNN751_2 1.368000
R3_110 Q_PNN751_3 Q_PNN751_4 4.000000
R4_110 Q_PNN751_5 Q_PNN751_4 0.304000
R5_110 Q_PNN751_5 Q_PNN751_6 4.000000
R6_110 Q_PNN751_7 Q_PNN751_6 0.304000
R7_110 Q_PNN751_7 U268:Z 4.000000

C1_40 iDFF_24_q_reg:Q 0 0.000045PF
C2_40 INP_PNN93_14 0 0.000105PF
C3_40 INP_PNN93_11 0 0.000105PF
C4_40 INP_PNN93_8 0 0.001035PF
C5_40 INP_PNN93_6 0 0.000984PF
C6_40 INP_PNN93_4 0 0.000121PF
C7_40 clk_r_REG43_S2:D 0 0.000045PF
C8_40 INP_PNN93_15 0 0.000044PF
C9_40 INP_PNN93_13 0 0.000044PF
C10_40 INP_PNN93_10 0 0.000069PF
C11_40 U213:A 0 0.000045PF
C12_40 INP_PNN93_9 0 0.000055PF
C13_40 INP_PNN93_7 0 0.000071PF
C14_40 INP_PNN93_5 0 0.000255PF
C15_40 INP_PNN93_3 0 0.000255PF
C16_40 INP_PNN93_2 0 0.000121PF
C17_40 U209:A 0 0.000090PF
R1_40 U209:A INP_PNN93_2 4.000000
R2_40 INP_PNN93_2 INP_PNN93_3 4.000000
R3_40 U209:A INP_PNN93_4 4.000000
R4_40 INP_PNN93_5 INP_PNN93_3 1.976000
R5_40 INP_PNN93_4 INP_PNN93_6 4.000000
R6_40 INP_PNN93_5 INP_PNN93_7 4.000000
R7_40 INP_PNN93_6 INP_PNN93_8 8.056000
R8_40 INP_PNN93_7 INP_PNN93_9 0.152000
R9_40 INP_PNN93_8 INP_PNN93_10 0.608000
R10_40 INP_PNN93_8 INP_PNN93_11 4.000000
R11_40 INP_PNN93_9 U213:A 4.000000
R12_40 INP_PNN93_10 INP_PNN93_13 4.000000
R13_40 INP_PNN93_11 INP_PNN93_14 1.064000
R14_40 INP_PNN93_15 INP_PNN93_13 0.304000
R15_40 INP_PNN93_14 iDFF_24_q_reg:Q 4.000000
R16_40 INP_PNN93_15 clk_r_REG43_S2:D 4.000000

C1_8 U200:B 0 0.000045PF
C2_8 INP_PNN121_8 0 0.000620PF
C3_8 INP_PNN121_11 0 0.000373PF
C4_8 INP_PNN121_14 0 0.000173PF
C5_8 INP_PNN121_15 0 0.000173PF
C6_8 INP_PNN121_16 0 0.000121PF
C7_8 U217:B 0 0.000045PF
C8_8 iDFF_31_q_reg:Q 0 0.000045PF
C9_8 INP_PNN121_10 0 0.000091PF
C10_8 INP_PNN121_7 0 0.000091PF
C11_8 INP_PNN121_4 0 0.000079PF
C12_8 INP_PNN121_2 0 0.000464PF
C13_8 INP_PNN121_5 0 0.000266PF
C14_8 clk_r_REG50_S2:D 0 0.000045PF
C15_8 INP_PNN121_6 0 0.000052PF
C16_8 INP_PNN121_3 0 0.000052PF
C17_8 INP_PNN121_1 0 0.000404PF
R1_8 INP_PNN121_1 INP_PNN121_2 3.952000
R2_8 INP_PNN121_1 INP_PNN121_3 4.000000
R3_8 INP_PNN121_2 INP_PNN121_4 0.608000
R4_8 INP_PNN121_2 INP_PNN121_5 4.000000
R5_8 INP_PNN121_6 INP_PNN121_3 0.456000
R6_8 INP_PNN121_4 INP_PNN121_7 4.000000
R7_8 INP_PNN121_8 INP_PNN121_5 2.736000
R8_8 INP_PNN121_6 clk_r_REG50_S2:D 4.000000
R9_8 INP_PNN121_7 INP_PNN121_10 0.912000
R10_8 INP_PNN121_11 INP_PNN121_8 1.824000
R11_8 INP_PNN121_8 U200:B 4.000000
R12_8 INP_PNN121_10 iDFF_31_q_reg:Q 4.000000
R13_8 INP_PNN121_11 INP_PNN121_14 4.000000
R14_8 INP_PNN121_14 INP_PNN121_15 1.520000
R15_8 INP_PNN121_15 INP_PNN121_16 4.000000
R16_8 INP_PNN121_16 U217:B 4.000000

C1_9 iDFF_32_q_reg:Q 0 0.000045PF
C2_9 INP_PNN125_14 0 0.000061PF
C3_9 INP_PNN125_11 0 0.000061PF
C4_9 INP_PNN125_8 0 0.000439PF
C5_9 INP_PNN125_5 0 0.000363PF
C6_9 INP_PNN125_2 0 0.000284PF
C7_9 INP_PNN125_4 0 0.000258PF
C8_9 U200:A 0 0.000045PF
C9_9 U207:B 0 0.000045PF
C10_9 INP_PNN125_16 0 0.000139PF
C11_9 INP_PNN125_13 0 0.000139PF
C12_9 INP_PNN125_10 0 0.000094PF
C13_9 clk_r_REG51_S2:D 0 0.000045PF
C14_9 INP_PNN125_12 0 0.000057PF
C15_9 INP_PNN125_9 0 0.000057PF
C16_9 INP_PNN125_6 0 0.000367PF
C17_9 INP_PNN125_3 0 0.000367PF
C18_9 INP_PNN125_1 0 0.000045PF
R1_9 INP_PNN125_2 INP_PNN125_1 0.304000
R2_9 INP_PNN125_1 INP_PNN125_3 4.000000
R3_9 INP_PNN125_4 INP_PNN125_2 2.584000
R4_9 INP_PNN125_2 INP_PNN125_5 4.000000
R5_9 INP_PNN125_6 INP_PNN125_3 3.800000
R6_9 INP_PNN125_4 U200:A 4.000000
R7_9 INP_PNN125_5 INP_PNN125_8 3.648000
R8_9 INP_PNN125_6 INP_PNN125_9 4.000000
R9_9 INP_PNN125_8 INP_PNN125_10 0.912000
R10_9 INP_PNN125_8 INP_PNN125_11 4.000000
R11_9 INP_PNN125_9 INP_PNN125_12 0.456000
R12_9 INP_PNN125_10 INP_PNN125_13 4.000000
R13_9 INP_PNN125_11 INP_PNN125_14 0.456000
R14_9 INP_PNN125_12 clk_r_REG51_S2:D 4.000000
R15_9 INP_PNN125_16 INP_PNN125_13 1.064000
R16_9 INP_PNN125_14 iDFF_32_q_reg:Q 4.000000
R17_9 INP_PNN125_16 U207:B 4.000000

C1_38 U213:B 0 0.000045PF
C2_38 INP_PNN89_8 0 0.000208PF
C3_38 INP_PNN89_10 0 0.000176PF
C4_38 INP_PNN89_13 0 0.000431PF
C5_38 INP_PNN89_15 0 0.000397PF
C6_38 U219:A 0 0.000045PF
C7_38 iDFF_23_q_reg:Q 0 0.000045PF
C8_38 INP_PNN89_12 0 0.000034PF
C9_38 INP_PNN89_9 0 0.000050PF
C10_38 INP_PNN89_7 0 0.000273PF
C11_38 INP_PNN89_5 0 0.000273PF
C12_38 INP_PNN89_2 0 0.000109PF
C13_38 INP_PNN89_4 0 0.000104PF
C14_38 INP_PNN89_6 0 0.000119PF
C15_38 clk_r_REG42_S2:D 0 0.000045PF
C16_38 INP_PNN89_1 0 0.000057PF
R1_38 INP_PNN89_2 INP_PNN89_1 0.456000
R2_38 INP_PNN89_1 clk_r_REG42_S2:D 4.000000
R3_38 INP_PNN89_4 INP_PNN89_2 0.608000
R4_38 INP_PNN89_2 INP_PNN89_5 4.000000
R5_38 INP_PNN89_6 INP_PNN89_4 0.152000
R6_38 INP_PNN89_5 INP_PNN89_7 2.128000
R7_38 INP_PNN89_8 INP_PNN89_6 0.912000
R8_38 INP_PNN89_7 INP_PNN89_9 4.000000
R9_38 INP_PNN89_10 INP_PNN89_8 1.520000
R10_38 INP_PNN89_8 U213:B 4.000000
R11_38 INP_PNN89_9 INP_PNN89_12 0.152000
R12_38 INP_PNN89_13 INP_PNN89_10 0.152000
R13_38 INP_PNN89_12 iDFF_23_q_reg:Q 4.000000
R14_38 INP_PNN89_15 INP_PNN89_13 1.824000
R15_38 INP_PNN89_15 U219:A 4.000000

C1_245 U278:A 0 0.000045PF
C2_245 n24_5 0 0.000121PF
C3_245 n24_4 0 0.000130PF
C4_245 n24_3 0 0.000130PF
C5_245 n24_2 0 0.000121PF
C6_245 clk_r_REG42_S2:Q 0 0.000045PF
R1_245 clk_r_REG42_S2:Q n24_2 4.000000
R2_245 n24_2 n24_3 4.000000
R3_245 n24_4 n24_3 1.976000
R4_245 n24_4 n24_5 4.000000
R5_245 n24_5 U278:A 4.000000

C1_311 U279:Z 0 0.000045PF
C2_311 n85_7 0 0.000444PF
C3_311 n85_6 0 0.000444PF
C4_311 n85_5 0 0.000057PF
C5_311 n85_4 0 0.000057PF
C6_311 n85_3 0 0.000071PF
C7_311 n85_2 0 0.000055PF
C8_311 U278:B 0 0.000045PF
R1_311 U278:B n85_2 4.000000
R2_311 n85_3 n85_2 0.152000
R3_311 n85_3 n85_4 4.000000
R4_311 n85_5 n85_4 0.456000
R5_311 n85_5 n85_6 4.000000
R6_311 n85_7 n85_6 3.800000
R7_311 n85_7 U279:Z 4.000000

C1_81 PNN93 0 0.001934PF
C2_81 PNN93_5 0 0.001990PF
C3_81 PNN93_4 0 0.000598PF
C4_81 PNN93_3 0 0.000563PF
C5_81 PNN93_2 0 0.000121PF
C6_81 iDFF_24_q_reg:D 0 0.000045PF
R1_81 iDFF_24_q_reg:D PNN93_2 4.000000
R2_81 PNN93_2 PNN93_3 4.000000
R3_81 PNN93_3 PNN93_4 7.144000
R4_81 PNN93_5 PNN93_4 0.152000
R5_81 PNN93_5 PNN93 24.471999

C1_105 U278:Z 0 0.000045PF
C2_105 Q_PNN746_7 0 0.000037PF
C3_105 Q_PNN746_6 0 0.000053PF
C4_105 Q_PNN746_5 0 0.000061PF
C5_105 Q_PNN746_4 0 0.000061PF
C6_105 Q_PNN746_3 0 0.000235PF
C7_105 Q_PNN746_2 0 0.000235PF
C8_105 oDFF_23_q_reg:D 0 0.000045PF
R1_105 oDFF_23_q_reg:D Q_PNN746_2 4.000000
R2_105 Q_PNN746_3 Q_PNN746_2 1.824000
R3_105 Q_PNN746_3 Q_PNN746_4 4.000000
R4_105 Q_PNN746_5 Q_PNN746_4 0.760000
R5_105 Q_PNN746_5 Q_PNN746_6 4.000000
R6_105 Q_PNN746_7 Q_PNN746_6 0.152000
R7_105 Q_PNN746_7 U278:Z 4.000000

C1_134 oDFF_20_q_reg:Q 0 0.000045PF
C2_134 Qout_PNN743_5 0 0.002424PF
C3_134 Qout_PNN743_4 0 0.002424PF
C4_134 Qout_PNN743_3 0 0.000044PF
C5_134 Qout_PNN743_2 0 0.000044PF
C6_134 Qout_PNN743 0 0.000042PF
R1_134 Qout_PNN743 Qout_PNN743_2 4.000000
R2_134 Qout_PNN743_3 Qout_PNN743_2 0.304000
R3_134 Qout_PNN743_3 Qout_PNN743_4 4.000000
R4_134 Qout_PNN743_5 Qout_PNN743_4 30.703999
R5_134 Qout_PNN743_5 oDFF_20_q_reg:Q 4.000000

C1_143 oDFF_29_q_reg:Q 0 0.000045PF
C2_143 Qout_PNN752_7 0 0.000044PF
C3_143 Qout_PNN752_6 0 0.000044PF
C4_143 Qout_PNN752_5 0 0.002494PF
C5_143 Qout_PNN752_4 0 0.002494PF
C6_143 Qout_PNN752_3 0 0.000044PF
C7_143 Qout_PNN752_2 0 0.000044PF
C8_143 Qout_PNN752 0 0.000042PF
R1_143 Qout_PNN752 Qout_PNN752_2 4.000000
R2_143 Qout_PNN752_2 Qout_PNN752_3 0.304000
R3_143 Qout_PNN752_3 Qout_PNN752_4 4.000000
R4_143 Qout_PNN752_4 Qout_PNN752_5 32.527999
R5_143 Qout_PNN752_5 Qout_PNN752_6 4.000000
R6_143 Qout_PNN752_7 Qout_PNN752_6 0.304000
R7_143 Qout_PNN752_7 oDFF_29_q_reg:Q 4.000000

C1_139 oDFF_25_q_reg:Q 0 0.000045PF
C2_139 Qout_PNN748_7 0 0.000039PF
C3_139 Qout_PNN748_6 0 0.000039PF
C4_139 Qout_PNN748_5 0 0.002364PF
C5_139 Qout_PNN748_4 0 0.002364PF
C6_139 Qout_PNN748_3 0 0.000044PF
C7_139 Qout_PNN748_2 0 0.000044PF
C8_139 Qout_PNN748 0 0.000042PF
R1_139 Qout_PNN748 Qout_PNN748_2 4.000000
R2_139 Qout_PNN748_2 Qout_PNN748_3 0.304000
R3_139 Qout_PNN748_3 Qout_PNN748_4 4.000000
R4_139 Qout_PNN748_4 Qout_PNN748_5 30.855999
R5_139 Qout_PNN748_5 Qout_PNN748_6 4.000000
R6_139 Qout_PNN748_7 Qout_PNN748_6 0.304000
R7_139 Qout_PNN748_7 oDFF_25_q_reg:Q 4.000000

C1_122 oDFF_8_q_reg:Q 0 0.000045PF
C2_122 Qout_PNN731_10 0 0.000121PF
C3_122 Qout_PNN731_9 0 0.000512PF
C4_122 Qout_PNN731_8 0 0.000512PF
C5_122 Qout_PNN731_7 0 0.000044PF
C6_122 Qout_PNN731_6 0 0.000044PF
C7_122 Qout_PNN731_5 0 0.002197PF
C8_122 Qout_PNN731_4 0 0.002197PF
C9_122 Qout_PNN731_3 0 0.000044PF
C10_122 Qout_PNN731_2 0 0.000044PF
C11_122 Qout_PNN731 0 0.000042PF
R1_122 Qout_PNN731 Qout_PNN731_2 4.000000
R2_122 Qout_PNN731_2 Qout_PNN731_3 0.304000
R3_122 Qout_PNN731_3 Qout_PNN731_4 4.000000
R4_122 Qout_PNN731_4 Qout_PNN731_5 27.815999
R5_122 Qout_PNN731_5 Qout_PNN731_6 4.000000
R6_122 Qout_PNN731_7 Qout_PNN731_6 0.304000
R7_122 Qout_PNN731_7 Qout_PNN731_8 4.000000
R8_122 Qout_PNN731_8 Qout_PNN731_9 5.624000
R9_122 Qout_PNN731_9 Qout_PNN731_10 4.000000
R10_122 Qout_PNN731_10 oDFF_8_q_reg:Q 4.000000

C1_42 PNN1 0 0.002315PF
C2_42 PNN1_8 0 0.002336PF
C3_42 PNN1_7 0 0.000045PF
C4_42 PNN1_6 0 0.000045PF
C5_42 PNN1_5 0 0.000690PF
C6_42 PNN1_4 0 0.000690PF
C7_42 PNN1_3 0 0.000051PF
C8_42 PNN1_2 0 0.000051PF
C9_42 iDFF_1_q_reg:D 0 0.000045PF
R1_42 iDFF_1_q_reg:D PNN1_2 4.000000
R2_42 PNN1_2 PNN1_3 0.304000
R3_42 PNN1_3 PNN1_4 4.000000
R4_42 PNN1_5 PNN1_4 6.840000
R5_42 PNN1_5 PNN1_6 4.000000
R6_42 PNN1_7 PNN1_6 0.304000
R7_42 PNN1_7 PNN1_8 4.000000
R8_42 PNN1 PNN1_8 28.727999

C1_299 U261:B 0 0.000045PF
C2_299 n74_26 0 0.000121PF
C3_299 n74_25 0 0.000394PF
C4_299 n74_23 0 0.000394PF
C5_299 n74_22 0 0.000108PF
C6_299 U263:B 0 0.000045PF
C7_299 U265:B 0 0.000045PF
C8_299 n74_2 0 0.000110PF
C9_299 n74_4 0 0.000121PF
C10_299 n74_7 0 0.000093PF
C11_299 n74_8 0 0.000093PF
C12_299 n74_9 0 0.000121PF
C13_299 n74_10 0 0.000763PF
C14_299 n74_11 0 0.000763PF
C15_299 n74_12 0 0.000197PF
C16_299 n74_13 0 0.000197PF
C17_299 n74_14 0 0.000057PF
C18_299 n74_15 0 0.000057PF
C19_299 U267:B 0 0.000090PF
C20_299 n74_17 0 0.000039PF
C21_299 n74_18 0 0.000055PF
C22_299 n74_19 0 0.000146PF
C23_299 n74_20 0 0.000146PF
C24_299 n74_21 0 0.000108PF
C25_299 U203:Z 0 0.000037PF
C26_299 n74_3 0 0.000060PF
C27_299 n74_1 0 0.000110PF
R1_299 n74_1 n74_2 0.912000
R2_299 n74_1 n74_3 4.000000
R3_299 n74_2 n74_4 4.000000
R4_299 n74_2 U265:B 4.000000
R5_299 U203:Z n74_3 0.304000
R6_299 n74_4 n74_7 4.000000
R7_299 n74_7 n74_8 0.912000
R8_299 n74_8 n74_9 4.000000
R9_299 n74_9 n74_10 4.000000
R10_299 n74_10 n74_11 5.320000
R11_299 n74_11 n74_12 4.000000
R12_299 n74_12 n74_13 0.912000
R13_299 n74_13 n74_14 4.000000
R14_299 n74_14 n74_15 0.456000
R15_299 n74_15 U267:B 4.000000
R16_299 U267:B n74_17 4.000000
R17_299 n74_17 n74_18 0.152000
R18_299 n74_18 n74_19 4.000000
R19_299 n74_19 n74_20 1.064000
R20_299 n74_20 n74_21 4.000000
R21_299 n74_21 n74_22 0.760000
R22_299 n74_22 n74_23 4.000000
R23_299 n74_22 U263:B 4.000000
R24_299 n74_23 n74_25 1.672000
R25_299 n74_25 n74_26 4.000000
R26_299 n74_26 U261:B 4.000000

C1_304 U271:B 0 0.000045PF
C2_304 n79_8 0 0.000121PF
C3_304 n79_4 0 0.000056PF
C4_304 n79_7 0 0.000090PF
C5_304 n79_11 0 0.000090PF
C6_304 n79_14 0 0.000587PF
C7_304 n79_16 0 0.000587PF
C8_304 n79_18 0 0.000050PF
C9_304 n79_20 0 0.000033PF
C10_304 U269:B 0 0.000045PF
C11_304 U273:B 0 0.000045PF
C12_304 n79_21 0 0.000097PF
C13_304 n79_19 0 0.000121PF
C14_304 n79_17 0 0.000093PF
C15_304 n79_15 0 0.000093PF
C16_304 n79_13 0 0.000121PF
C17_304 n79_9 0 0.000861PF
C18_304 n79_5 0 0.000861PF
C19_304 n79_2 0 0.000203PF
C20_304 U204:Z 0 0.000045PF
C21_304 n79_27 0 0.000121PF
C22_304 n79_26 0 0.000096PF
C23_304 n79_25 0 0.000096PF
C24_304 n79_23 0 0.000097PF
C25_304 U275:B 0 0.000045PF
C26_304 n79_6 0 0.000143PF
C27_304 n79_3 0 0.000143PF
C28_304 n79_1 0 0.000166PF
R1_304 n79_1 n79_2 1.368000
R2_304 n79_1 n79_3 4.000000
R3_304 n79_2 n79_4 0.304000
R4_304 n79_2 n79_5 4.000000
R5_304 n79_3 n79_6 1.064000
R6_304 n79_4 n79_7 4.000000
R7_304 n79_4 n79_8 4.000000
R8_304 n79_9 n79_5 5.928000
R9_304 n79_6 U275:B 4.000000
R10_304 n79_7 n79_11 0.912000
R11_304 n79_8 U271:B 4.000000
R12_304 n79_9 n79_13 4.000000
R13_304 n79_11 n79_14 4.000000
R14_304 n79_13 n79_15 4.000000
R15_304 n79_14 n79_16 3.648000
R16_304 n79_17 n79_15 0.912000
R17_304 n79_16 n79_18 4.000000
R18_304 n79_17 n79_19 4.000000
R19_304 n79_18 n79_20 0.152000
R20_304 n79_19 n79_21 4.000000
R21_304 n79_20 U269:B 4.000000
R22_304 n79_23 n79_21 0.912000
R23_304 n79_21 U273:B 4.000000
R24_304 n79_23 n79_25 4.000000
R25_304 n79_26 n79_25 0.760000
R26_304 n79_26 n79_27 4.000000
R27_304 n79_27 U204:Z 4.000000

C1_7 U257:B 0 0.000045PF
C2_7 INP_PNN117_19 0 0.000121PF
C3_7 INP_PNN117_18 0 0.000287PF
C4_7 INP_PNN117_16 0 0.000287PF
C5_7 INP_PNN117_15 0 0.000128PF
C6_7 U199:B 0 0.000045PF
C7_7 clk_r_REG49_S2:D 0 0.000045PF
C8_7 INP_PNN117_8 0 0.000049PF
C9_7 INP_PNN117_5 0 0.000049PF
C10_7 INP_PNN117_2 0 0.000749PF
C11_7 INP_PNN117_4 0 0.000230PF
C12_7 INP_PNN117_7 0 0.000046PF
C13_7 INP_PNN117_10 0 0.000046PF
C14_7 INP_PNN117_12 0 0.001265PF
C15_7 INP_PNN117_13 0 0.001265PF
C16_7 INP_PNN117_14 0 0.000112PF
C17_7 iDFF_30_q_reg:Q 0 0.000045PF
C18_7 INP_PNN117_6 0 0.000054PF
C19_7 INP_PNN117_3 0 0.000071PF
C20_7 INP_PNN117_1 0 0.000538PF
R1_7 INP_PNN117_1 INP_PNN117_2 2.584000
R2_7 INP_PNN117_1 INP_PNN117_3 4.000000
R3_7 INP_PNN117_2 INP_PNN117_4 1.976000
R4_7 INP_PNN117_2 INP_PNN117_5 4.000000
R5_7 INP_PNN117_6 INP_PNN117_3 0.152000
R6_7 INP_PNN117_4 INP_PNN117_7 4.000000
R7_7 INP_PNN117_8 INP_PNN117_5 0.304000
R8_7 INP_PNN117_6 iDFF_30_q_reg:Q 4.000000
R9_7 INP_PNN117_7 INP_PNN117_10 0.304000
R10_7 INP_PNN117_8 clk_r_REG49_S2:D 4.000000
R11_7 INP_PNN117_10 INP_PNN117_12 4.000000
R12_7 INP_PNN117_12 INP_PNN117_13 10.336000
R13_7 INP_PNN117_13 INP_PNN117_14 4.000000
R14_7 INP_PNN117_15 INP_PNN117_14 0.912000
R15_7 INP_PNN117_15 INP_PNN117_16 4.000000
R16_7 INP_PNN117_15 U199:B 4.000000
R17_7 INP_PNN117_16 INP_PNN117_18 2.584000
R18_7 INP_PNN117_18 INP_PNN117_19 4.000000
R19_7 INP_PNN117_19 U257:B 4.000000

C1_141 oDFF_27_q_reg:Q 0 0.000045PF
C2_141 Qout_PNN750_11 0 0.000214PF
C3_141 Qout_PNN750_10 0 0.000214PF
C4_141 Qout_PNN750_9 0 0.000121PF
C5_141 Qout_PNN750_8 0 0.000063PF
C6_141 Qout_PNN750_7 0 0.000063PF
C7_141 Qout_PNN750_6 0 0.000121PF
C8_141 Qout_PNN750_5 0 0.002705PF
C9_141 Qout_PNN750_4 0 0.002705PF
C10_141 Qout_PNN750_3 0 0.000046PF
C11_141 Qout_PNN750_2 0 0.000046PF
C12_141 Qout_PNN750 0 0.000042PF
R1_141 Qout_PNN750 Qout_PNN750_2 4.000000
R2_141 Qout_PNN750_3 Qout_PNN750_2 0.304000
R3_141 Qout_PNN750_3 Qout_PNN750_4 4.000000
R4_141 Qout_PNN750_5 Qout_PNN750_4 33.135999
R5_141 Qout_PNN750_5 Qout_PNN750_6 4.000000
R6_141 Qout_PNN750_6 Qout_PNN750_7 4.000000
R7_141 Qout_PNN750_8 Qout_PNN750_7 0.608000
R8_141 Qout_PNN750_8 Qout_PNN750_9 4.000000
R9_141 Qout_PNN750_9 Qout_PNN750_10 4.000000
R10_141 Qout_PNN750_11 Qout_PNN750_10 2.888000
R11_141 Qout_PNN750_11 oDFF_27_q_reg:Q 4.000000

C1_175 U230:B 0 0.000045PF
C2_175 n110_20 0 0.000086PF
C3_175 n110_17 0 0.000436PF
C4_175 n110_15 0 0.000235PF
C5_175 n110_13 0 0.002154PF
C6_175 n110_11 0 0.002154PF
C7_175 n110_9 0 0.000496PF
C8_175 n110_7 0 0.000126PF
C9_175 n110_4 0 0.000752PF
C10_175 n110_2 0 0.001283PF
C11_175 n110_5 0 0.000121PF
C12_175 U247:B 0 0.000045PF
C13_175 U233:B 0 0.000045PF
C14_175 n110_19 0 0.000188PF
C15_175 U163:Z 0 0.000045PF
C16_175 n110_16 0 0.000121PF
C17_175 n110_14 0 0.000039PF
C18_175 n110_12 0 0.000055PF
C19_175 n110_10 0 0.000389PF
C20_175 U241:B 0 0.000045PF
C21_175 n110_3 0 0.000121PF
C22_175 n110_1 0 0.000550PF
R1_175 n110_1 n110_2 2.584000
R2_175 n110_1 n110_3 4.000000
R3_175 n110_2 n110_4 2.584000
R4_175 n110_2 n110_5 4.000000
R5_175 n110_3 U241:B 4.000000
R6_175 n110_4 n110_7 4.000000
R7_175 n110_5 U247:B 4.000000
R8_175 n110_7 n110_9 1.216000
R9_175 n110_9 n110_10 4.712000
R10_175 n110_9 n110_11 4.000000
R11_175 n110_10 n110_12 4.000000
R12_175 n110_11 n110_13 19.759999
R13_175 n110_12 n110_14 0.152000
R14_175 n110_13 n110_15 4.000000
R15_175 n110_14 n110_16 4.000000
R16_175 n110_17 n110_15 1.368000
R17_175 n110_16 U163:Z 4.000000
R18_175 n110_19 n110_17 1.064000
R19_175 n110_17 n110_20 0.152000
R20_175 n110_19 U233:B 4.000000
R21_175 n110_20 U230:B 4.000000

C1_68 PNN49 0 0.000042PF
C2_68 PNN49_7 0 0.000121PF
C3_68 PNN49_6 0 0.000538PF
C4_68 PNN49_5 0 0.000538PF
C5_68 PNN49_4 0 0.000121PF
C6_68 PNN49_3 0 0.002116PF
C7_68 PNN49_2 0 0.002116PF
C8_68 iDFF_13_q_reg:D 0 0.000045PF
R1_68 iDFF_13_q_reg:D PNN49_2 4.000000
R2_68 PNN49_3 PNN49_2 26.447999
R3_68 PNN49_3 PNN49_4 4.000000
R4_68 PNN49_4 PNN49_5 4.000000
R5_68 PNN49_6 PNN49_5 6.536000
R6_68 PNN49_6 PNN49_7 4.000000
R7_68 PNN49_7 PNN49 4.000000

C1_142 oDFF_28_q_reg:Q 0 0.000045PF
C2_142 Qout_PNN751_8 0 0.002131PF
C3_142 Qout_PNN751_7 0 0.002131PF
C4_142 Qout_PNN751_6 0 0.000121PF
C5_142 Qout_PNN751_5 0 0.000574PF
C6_142 Qout_PNN751_4 0 0.000574PF
C7_142 Qout_PNN751_3 0 0.000044PF
C8_142 Qout_PNN751_2 0 0.000044PF
C9_142 Qout_PNN751 0 0.000042PF
R1_142 Qout_PNN751 Qout_PNN751_2 4.000000
R2_142 Qout_PNN751_3 Qout_PNN751_2 0.304000
R3_142 Qout_PNN751_3 Qout_PNN751_4 4.000000
R4_142 Qout_PNN751_5 Qout_PNN751_4 6.992000
R5_142 Qout_PNN751_5 Qout_PNN751_6 4.000000
R6_142 Qout_PNN751_6 Qout_PNN751_7 4.000000
R7_142 Qout_PNN751_8 Qout_PNN751_7 25.687999
R8_142 Qout_PNN751_8 oDFF_28_q_reg:Q 4.000000

C1_158 U169:A 0 0.000045PF
C2_158 c0_n52_26 0 0.000064PF
C3_158 c0_n52_24 0 0.000064PF
C4_158 c0_n52_22 0 0.000405PF
C5_158 c0_n52_21 0 0.000323PF
C6_158 c0_n52_20 0 0.000177PF
C7_158 c0_n52_19 0 0.000177PF
C8_158 c0_n52_18 0 0.001928PF
C9_158 c0_n52_16 0 0.001928PF
C10_158 c0_n52_14 0 0.000253PF
C11_158 c0_n52_15 0 0.000161PF
C12_158 clk_r_REG20_S2:D 0 0.000045PF
C13_158 U189:B 0 0.000045PF
C14_158 c0_n52_36 0 0.000283PF
C15_158 c0_n52_35 0 0.000283PF
C16_158 c0_n52_34 0 0.000375PF
C17_158 c0_n52_33 0 0.000375PF
C18_158 c0_n52_32 0 0.000121PF
C19_158 U185:A 0 0.000090PF
C20_158 c0_n52_30 0 0.000215PF
C21_158 c0_n52_29 0 0.000215PF
C22_158 c0_n52_27 0 0.000763PF
C23_158 c0_n52_25 0 0.000797PF
C24_158 c0_n52_23 0 0.000136PF
C25_158 U243:A 0 0.000045PF
C26_158 c0_n52_3 0 0.000379PF
C27_158 c0_n52_5 0 0.000317PF
C28_158 U230:A 0 0.000090PF
C29_158 c0_n52_9 0 0.000121PF
C30_158 c0_n52_10 0 0.000121PF
C31_158 c0_n52_11 0 0.000090PF
C32_158 c0_n52_12 0 0.000090PF
C33_158 c0_n52_13 0 0.000110PF
C34_158 U159:Z 0 0.000045PF
C35_158 c0_n52_4 0 0.000121PF
C36_158 c0_n52_2 0 0.000440PF
C37_158 c0_n52_1 0 0.000440PF
R1_158 c0_n52_2 c0_n52_1 2.736000
R2_158 c0_n52_1 c0_n52_3 4.000000
R3_158 c0_n52_2 c0_n52_4 4.000000
R4_158 c0_n52_5 c0_n52_3 2.432000
R5_158 c0_n52_3 U243:A 4.000000
R6_158 c0_n52_4 U159:Z 4.000000
R7_158 c0_n52_5 U230:A 4.000000
R8_158 U230:A c0_n52_9 4.000000
R9_158 c0_n52_10 c0_n52_9 0.456000
R10_158 c0_n52_10 c0_n52_11 4.000000
R11_158 c0_n52_12 c0_n52_11 0.304000
R12_158 c0_n52_12 c0_n52_13 4.000000
R13_158 c0_n52_14 c0_n52_13 1.672000
R14_158 c0_n52_15 c0_n52_14 1.520000
R15_158 c0_n52_14 c0_n52_16 4.000000
R16_158 c0_n52_15 clk_r_REG20_S2:D 4.000000
R17_158 c0_n52_18 c0_n52_16 17.935999
R18_158 c0_n52_18 c0_n52_19 4.000000
R19_158 c0_n52_19 c0_n52_20 1.976000
R20_158 c0_n52_20 c0_n52_21 4.000000
R21_158 c0_n52_22 c0_n52_21 1.368000
R22_158 c0_n52_23 c0_n52_22 0.608000
R23_158 c0_n52_22 c0_n52_24 4.000000
R24_158 c0_n52_23 c0_n52_25 0.152000
R25_158 c0_n52_24 c0_n52_26 0.456000
R26_158 c0_n52_27 c0_n52_25 3.344000
R27_158 c0_n52_26 U169:A 4.000000
R28_158 c0_n52_27 c0_n52_29 4.000000
R29_158 c0_n52_29 c0_n52_30 2.280000
R30_158 c0_n52_30 U185:A 4.000000
R31_158 U185:A c0_n52_32 4.000000
R32_158 c0_n52_32 c0_n52_33 4.000000
R33_158 c0_n52_34 c0_n52_33 1.672000
R34_158 c0_n52_34 c0_n52_35 4.000000
R35_158 c0_n52_35 c0_n52_36 1.520000
R36_158 c0_n52_36 U189:B 4.000000

C1_285 U166:C 0 0.000045PF
C2_285 n61_13 0 0.000260PF
C3_285 n61_15 0 0.000216PF
C4_285 n61_17 0 0.000121PF
C5_285 n61_18 0 0.000104PF
C6_285 n61_19 0 0.000104PF
C7_285 n61_20 0 0.000320PF
C8_285 n61_21 0 0.000320PF
C9_285 n61_22 0 0.000135PF
C10_285 n61_23 0 0.000135PF
C11_285 U162:C 0 0.000045PF
C12_285 U168:C 0 0.000045PF
C13_285 n61_12 0 0.000491PF
C14_285 n61_8 0 0.000491PF
C15_285 n61_4 0 0.000486PF
C16_285 n61_7 0 0.000416PF
C17_285 n61_11 0 0.000063PF
C18_285 U181:Z 0 0.000045PF
C19_285 n61_5 0 0.000121PF
C20_285 n61_2 0 0.003023PF
C21_285 clk_r_REG28_S2:D 0 0.000045PF
C22_285 n61_6 0 0.000122PF
C23_285 n61_3 0 0.000122PF
C24_285 n61_1 0 0.002953PF
R1_285 n61_2 n61_1 14.896000
R2_285 n61_1 n61_3 4.000000
R3_285 n61_4 n61_2 0.304000
R4_285 n61_2 n61_5 4.000000
R5_285 n61_6 n61_3 1.976000
R6_285 n61_7 n61_4 1.824000
R7_285 n61_4 n61_8 4.000000
R8_285 n61_5 U181:Z 4.000000
R9_285 n61_6 clk_r_REG28_S2:D 4.000000
R10_285 n61_7 n61_11 4.000000
R11_285 n61_8 n61_12 3.648000
R12_285 n61_13 n61_11 0.304000
R13_285 n61_12 U168:C 4.000000
R14_285 n61_15 n61_13 0.760000
R15_285 n61_13 U166:C 4.000000
R16_285 n61_15 n61_17 4.000000
R17_285 n61_17 n61_18 4.000000
R18_285 n61_19 n61_18 1.520000
R19_285 n61_19 n61_20 4.000000
R20_285 n61_21 n61_20 3.040000
R21_285 n61_21 n61_22 4.000000
R22_285 n61_23 n61_22 1.976000
R23_285 n61_23 U162:C 4.000000

C1_130 oDFF_16_q_reg:Q 0 0.000045PF
C2_130 Qout_PNN739_8 0 0.000159PF
C3_130 Qout_PNN739_7 0 0.000159PF
C4_130 Qout_PNN739_6 0 0.000121PF
C5_130 Qout_PNN739_5 0 0.002266PF
C6_130 Qout_PNN739_4 0 0.002266PF
C7_130 Qout_PNN739_3 0 0.000113PF
C8_130 Qout_PNN739_2 0 0.000113PF
C9_130 Qout_PNN739 0 0.000042PF
R1_130 Qout_PNN739 Qout_PNN739_2 4.000000
R2_130 Qout_PNN739_3 Qout_PNN739_2 1.216000
R3_130 Qout_PNN739_3 Qout_PNN739_4 4.000000
R4_130 Qout_PNN739_4 Qout_PNN739_5 29.031999
R5_130 Qout_PNN739_5 Qout_PNN739_6 4.000000
R6_130 Qout_PNN739_6 Qout_PNN739_7 4.000000
R7_130 Qout_PNN739_7 Qout_PNN739_8 1.672000
R8_130 Qout_PNN739_8 oDFF_16_q_reg:Q 4.000000

C1_48 PNN121 0 0.002424PF
C2_48 PNN121_5 0 0.002445PF
C3_48 PNN121_4 0 0.000121PF
C4_48 PNN121_3 0 0.000632PF
C5_48 PNN121_2 0 0.000632PF
C6_48 iDFF_31_q_reg:D 0 0.000045PF
R1_48 iDFF_31_q_reg:D PNN121_2 4.000000
R2_48 PNN121_2 PNN121_3 2.736000
R3_48 PNN121_3 PNN121_4 4.000000
R4_48 PNN121_4 PNN121_5 4.000000
R5_48 PNN121_5 PNN121 30.399999

C1_50 PNN129 0 0.000042PF
C2_50 PNN129_13 0 0.000121PF
C3_50 PNN129_12 0 0.000573PF
C4_50 PNN129_11 0 0.000573PF
C5_50 PNN129_10 0 0.000121PF
C6_50 PNN129_9 0 0.002614PF
C7_50 PNN129_8 0 0.002614PF
C8_50 PNN129_7 0 0.000121PF
C9_50 PNN129_6 0 0.000605PF
C10_50 PNN129_5 0 0.000605PF
C11_50 PNN129_4 0 0.000121PF
C12_50 PNN129_3 0 0.000271PF
C13_50 PNN129_2 0 0.000271PF
C14_50 iDFF_33_q_reg:D 0 0.000045PF
R1_50 iDFF_33_q_reg:D PNN129_2 4.000000
R2_50 PNN129_3 PNN129_2 3.040000
R3_50 PNN129_3 PNN129_4 4.000000
R4_50 PNN129_4 PNN129_5 4.000000
R5_50 PNN129_6 PNN129_5 7.144000
R6_50 PNN129_6 PNN129_7 4.000000
R7_50 PNN129_7 PNN129_8 4.000000
R8_50 PNN129_9 PNN129_8 30.399999
R9_50 PNN129_9 PNN129_10 4.000000
R10_50 PNN129_10 PNN129_11 4.000000
R11_50 PNN129_12 PNN129_11 6.536000
R12_50 PNN129_12 PNN129_13 4.000000
R13_50 PNN129_13 PNN129 4.000000

C1_193 U180:B 0 0.000045PF
C2_193 n127_10 0 0.000264PF
C3_193 n127_8 0 0.000423PF
C4_193 n127_5 0 0.000423PF
C5_193 n127_2 0 0.000170PF
C6_193 n127_4 0 0.000048PF
C7_193 U176:B 0 0.000045PF
C8_193 U174:B 0 0.000045PF
C9_193 n127_19 0 0.000121PF
C10_193 n127_17 0 0.000078PF
C11_193 n127_15 0 0.000078PF
C12_193 n127_12 0 0.000201PF
C13_193 U199:Z 0 0.000045PF
C14_193 n127_18 0 0.000092PF
C15_193 n127_16 0 0.000092PF
C16_193 n127_14 0 0.000121PF
C17_193 n127_11 0 0.000503PF
C18_193 n127_9 0 0.000503PF
C19_193 n127_6 0 0.000133PF
C20_193 n127_3 0 0.000133PF
C21_193 n127_1 0 0.000141PF
R1_193 n127_2 n127_1 1.368000
R2_193 n127_1 n127_3 4.000000
R3_193 n127_4 n127_2 0.304000
R4_193 n127_2 n127_5 4.000000
R5_193 n127_6 n127_3 1.064000
R6_193 n127_4 U176:B 4.000000
R7_193 n127_5 n127_8 5.776000
R8_193 n127_6 n127_9 4.000000
R9_193 n127_8 n127_10 4.000000
R10_193 n127_9 n127_11 6.384000
R11_193 n127_12 n127_10 2.128000
R12_193 n127_10 U180:B 4.000000
R13_193 n127_11 n127_14 4.000000
R14_193 n127_12 n127_15 4.000000
R15_193 n127_14 n127_16 4.000000
R16_193 n127_15 n127_17 0.456000
R17_193 n127_16 n127_18 1.368000
R18_193 n127_17 n127_19 4.000000
R19_193 n127_18 U199:Z 4.000000
R20_193 n127_19 U174:B 4.000000

C1_168 U235:B 0 0.000093PF
C2_168 n104_5 0 0.000115PF
C3_168 n104_2 0 0.001144PF
C4_168 n104_4 0 0.000102PF
C5_168 U316:B 0 0.000045PF
C6_168 U243:B 0 0.000045PF
C7_168 n104_32 0 0.000293PF
C8_168 n104_31 0 0.000293PF
C9_168 n104_30 0 0.000957PF
C10_168 n104_29 0 0.000957PF
C11_168 n104_28 0 0.000117PF
C12_168 n104_27 0 0.000054PF
C13_168 U245:B 0 0.000090PF
C14_168 n104_25 0 0.000121PF
C15_168 n104_24 0 0.000401PF
C16_168 n104_23 0 0.000436PF
C17_168 n104_22 0 0.001028PF
C18_168 n104_21 0 0.000993PF
C19_168 n104_20 0 0.000064PF
C20_168 n104_19 0 0.000064PF
C21_168 n104_18 0 0.000368PF
C22_168 n104_17 0 0.000368PF
C23_168 n104_16 0 0.000075PF
C24_168 n104_15 0 0.000075PF
C25_168 n104_14 0 0.000497PF
C26_168 n104_13 0 0.000497PF
C27_168 n104_12 0 0.000077PF
C28_168 n104_11 0 0.000060PF
C29_168 U161:Z 0 0.000090PF
C30_168 n104_9 0 0.000121PF
C31_168 n104_6 0 0.000290PF
C32_168 n104_3 0 0.000290PF
C33_168 n104_1 0 0.001060PF
R1_168 n104_2 n104_1 10.184000
R2_168 n104_1 n104_3 4.000000
R3_168 n104_4 n104_2 0.912000
R4_168 n104_2 n104_5 4.000000
R5_168 n104_3 n104_6 3.800000
R6_168 n104_4 U316:B 4.000000
R7_168 U235:B n104_5 0.760000
R8_168 n104_6 n104_9 4.000000
R9_168 n104_9 U161:Z 4.000000
R10_168 U161:Z n104_11 4.000000
R11_168 n104_12 n104_11 0.152000
R12_168 n104_12 n104_13 4.000000
R13_168 n104_13 n104_14 4.408000
R14_168 n104_14 n104_15 4.000000
R15_168 n104_15 n104_16 0.456000
R16_168 n104_16 n104_17 4.000000
R17_168 n104_17 n104_18 2.280000
R18_168 n104_18 n104_19 4.000000
R19_168 n104_20 n104_19 0.456000
R20_168 n104_20 n104_21 4.000000
R21_168 n104_21 n104_22 8.208000
R22_168 n104_22 n104_23 0.152000
R23_168 n104_23 n104_24 2.432000
R24_168 n104_24 n104_25 4.000000
R25_168 n104_25 U245:B 4.000000
R26_168 U245:B n104_27 4.000000
R27_168 n104_28 n104_27 0.152000
R28_168 n104_28 n104_29 4.000000
R29_168 n104_29 n104_30 3.344000
R30_168 n104_30 n104_31 4.000000
R31_168 n104_32 n104_31 3.496000
R32_168 n104_32 U243:B 4.000000

C1_45 PNN109 0 0.002448PF
C2_45 PNN109_10 0 0.002469PF
C3_45 PNN109_9 0 0.000033PF
C4_45 PNN109_8 0 0.000049PF
C5_45 PNN109_7 0 0.000343PF
C6_45 PNN109_6 0 0.000343PF
C7_45 PNN109_5 0 0.000060PF
C8_45 PNN109_4 0 0.000044PF
C9_45 PNN109_3 0 0.000081PF
C10_45 PNN109_2 0 0.000081PF
C11_45 iDFF_28_q_reg:D 0 0.000045PF
R1_45 iDFF_28_q_reg:D PNN109_2 4.000000
R2_45 PNN109_2 PNN109_3 1.216000
R3_45 PNN109_3 PNN109_4 4.000000
R4_45 PNN109_5 PNN109_4 0.152000
R5_45 PNN109_5 PNN109_6 4.000000
R6_45 PNN109_6 PNN109_7 3.496000
R7_45 PNN109_7 PNN109_8 4.000000
R8_45 PNN109_8 PNN109_9 0.152000
R9_45 PNN109_9 PNN109_10 4.000000
R10_45 PNN109_10 PNN109 30.095999

C1_67 PNN45 0 0.000042PF
C2_67 PNN45_7 0 0.000121PF
C3_67 PNN45_6 0 0.000586PF
C4_67 PNN45_5 0 0.000586PF
C5_67 PNN45_4 0 0.000121PF
C6_67 PNN45_3 0 0.002622PF
C7_67 PNN45_2 0 0.002622PF
C8_67 iDFF_12_q_reg:D 0 0.000045PF
R1_67 iDFF_12_q_reg:D PNN45_2 4.000000
R2_67 PNN45_3 PNN45_2 30.247999
R3_67 PNN45_3 PNN45_4 4.000000
R4_67 PNN45_4 PNN45_5 4.000000
R5_67 PNN45_6 PNN45_5 6.688000
R6_67 PNN45_6 PNN45_7 4.000000
R7_67 PNN45_7 PNN45 4.000000

C1_49 PNN125 0 0.002512PF
C2_49 PNN125_5 0 0.002533PF
C3_49 PNN125_4 0 0.000121PF
C4_49 PNN125_3 0 0.000246PF
C5_49 PNN125_2 0 0.000246PF
C6_49 iDFF_32_q_reg:D 0 0.000045PF
R1_49 iDFF_32_q_reg:D PNN125_2 4.000000
R2_49 PNN125_2 PNN125_3 2.736000
R3_49 PNN125_3 PNN125_4 4.000000
R4_49 PNN125_4 PNN125_5 4.000000
R5_49 PNN125_5 PNN125 30.399999

C1_321 U295:B 0 0.000045PF
C2_321 n94_26 0 0.000121PF
C3_321 n94_25 0 0.000128PF
C4_321 n94_24 0 0.000128PF
C5_321 n94_23 0 0.000121PF
C6_321 U297:B 0 0.000090PF
C7_321 n94_21 0 0.000163PF
C8_321 n94_19 0 0.000163PF
C9_321 n94_17 0 0.001073PF
C10_321 n94_15 0 0.001073PF
C11_321 n94_12 0 0.000389PF
C12_321 n94_8 0 0.000389PF
C13_321 n94_5 0 0.000676PF
C14_321 n94_9 0 0.000121PF
C15_321 U293:B 0 0.000045PF
C16_321 U299:B 0 0.000045PF
C17_321 n94_6 0 0.000121PF
C18_321 n94_3 0 0.000676PF
C19_321 U210:Z 0 0.000045PF
C20_321 n94_18 0 0.000362PF
C21_321 n94_16 0 0.000396PF
C22_321 n94_14 0 0.001034PF
C23_321 n94_11 0 0.001000PF
C24_321 n94_7 0 0.000035PF
C25_321 n94_4 0 0.000051PF
C26_321 n94_2 0 0.000096PF
C27_321 n94_1 0 0.000096PF
R1_321 n94_1 n94_2 1.672000
R2_321 n94_1 n94_3 4.000000
R3_321 n94_2 n94_4 4.000000
R4_321 n94_3 n94_5 8.208000
R5_321 n94_3 n94_6 4.000000
R6_321 n94_7 n94_4 0.152000
R7_321 n94_5 n94_8 4.000000
R8_321 n94_5 n94_9 4.000000
R9_321 n94_6 U299:B 4.000000
R10_321 n94_7 n94_11 4.000000
R11_321 n94_8 n94_12 1.672000
R12_321 n94_9 U293:B 4.000000
R13_321 n94_11 n94_14 7.752000
R14_321 n94_12 n94_15 4.000000
R15_321 n94_16 n94_14 0.152000
R16_321 n94_15 n94_17 10.792000
R17_321 n94_16 n94_18 2.280000
R18_321 n94_17 n94_19 4.000000
R19_321 n94_18 U210:Z 4.000000
R20_321 n94_19 n94_21 0.912000
R21_321 n94_21 U297:B 4.000000
R22_321 U297:B n94_23 4.000000
R23_321 n94_23 n94_24 4.000000
R24_321 n94_24 n94_25 0.912000
R25_321 n94_25 n94_26 4.000000
R26_321 n94_26 U295:B 4.000000

C1_31 U253:A 0 0.000019PF
C2_31 INP_PNN61_20 0 0.000051PF
C3_31 INP_PNN61_18 0 0.000054PF
C4_31 INP_PNN61_16 0 0.000071PF
C5_31 INP_PNN61_14 0 0.000660PF
C6_31 INP_PNN61_11 0 0.000660PF
C7_31 INP_PNN61_8 0 0.000729PF
C8_31 INP_PNN61_10 0 0.000137PF
C9_31 INP_PNN61_13 0 0.000121PF
C10_31 INP_PNN61_15 0 0.000110PF
C11_31 INP_PNN61_17 0 0.000110PF
C12_31 U193:A 0 0.000045PF
C13_31 iDFF_16_q_reg:Q 0 0.000045PF
C14_31 INP_PNN61_9 0 0.000034PF
C15_31 INP_PNN61_7 0 0.000050PF
C16_31 INP_PNN61_4 0 0.000105PF
C17_31 INP_PNN61_2 0 0.000251PF
C18_31 INP_PNN61_5 0 0.000611PF
C19_31 clk_r_REG35_S2:D 0 0.000045PF
C20_31 INP_PNN61_3 0 0.000121PF
C21_31 INP_PNN61_1 0 0.000165PF
R1_31 INP_PNN61_1 INP_PNN61_2 1.064000
R2_31 INP_PNN61_1 INP_PNN61_3 4.000000
R3_31 INP_PNN61_2 INP_PNN61_4 1.064000
R4_31 INP_PNN61_2 INP_PNN61_5 4.000000
R5_31 INP_PNN61_3 clk_r_REG35_S2:D 4.000000
R6_31 INP_PNN61_4 INP_PNN61_7 4.000000
R7_31 INP_PNN61_5 INP_PNN61_8 4.408000
R8_31 INP_PNN61_7 INP_PNN61_9 0.152000
R9_31 INP_PNN61_8 INP_PNN61_10 1.824000
R10_31 INP_PNN61_8 INP_PNN61_11 4.000000
R11_31 INP_PNN61_9 iDFF_16_q_reg:Q 4.000000
R12_31 INP_PNN61_10 INP_PNN61_13 4.000000
R13_31 INP_PNN61_11 INP_PNN61_14 4.408000
R14_31 INP_PNN61_13 INP_PNN61_15 4.000000
R15_31 INP_PNN61_14 INP_PNN61_16 4.000000
R16_31 INP_PNN61_15 INP_PNN61_17 0.912000
R17_31 INP_PNN61_18 INP_PNN61_16 0.152000
R18_31 INP_PNN61_17 U193:A 4.000000
R19_31 INP_PNN61_18 INP_PNN61_20 4.000000
R20_31 INP_PNN61_20 U253:A 0.152000

C1_46 PNN113 0 0.000042PF
C2_46 PNN113_13 0 0.000121PF
C3_46 PNN113_12 0 0.000663PF
C4_46 PNN113_11 0 0.000663PF
C5_46 PNN113_10 0 0.000121PF
C6_46 PNN113_9 0 0.002292PF
C7_46 PNN113_8 0 0.002292PF
C8_46 PNN113_7 0 0.000121PF
C9_46 PNN113_6 0 0.000066PF
C10_46 PNN113_5 0 0.000066PF
C11_46 PNN113_4 0 0.000121PF
C12_46 PNN113_3 0 0.000948PF
C13_46 PNN113_2 0 0.000948PF
C14_46 iDFF_29_q_reg:D 0 0.000045PF
R1_46 iDFF_29_q_reg:D PNN113_2 4.000000
R2_46 PNN113_2 PNN113_3 7.296000
R3_46 PNN113_3 PNN113_4 4.000000
R4_46 PNN113_4 PNN113_5 4.000000
R5_46 PNN113_5 PNN113_6 0.760000
R6_46 PNN113_6 PNN113_7 4.000000
R7_46 PNN113_7 PNN113_8 4.000000
R8_46 PNN113_8 PNN113_9 27.055999
R9_46 PNN113_9 PNN113_10 4.000000
R10_46 PNN113_10 PNN113_11 4.000000
R11_46 PNN113_11 PNN113_12 7.600000
R12_46 PNN113_12 PNN113_13 4.000000
R13_46 PNN113_13 PNN113 4.000000

C1_161 clk 0 0.000042PF
C2_161 clk_7 0 0.000121PF
C3_161 clk_6 0 0.003609PF
C4_161 clk_5 0 0.003609PF
C5_161 clk_4 0 0.000511PF
C6_161 clk_3 0 0.000511PF
C7_161 clk_2 0 0.000121PF
C8_161 clk__L1_I0:A 0 0.000045PF
R1_161 clk__L1_I0:A clk_2 4.000000
R2_161 clk_2 clk_3 4.000000
R3_161 clk_4 clk_3 7.448000
R4_161 clk_4 clk_5 4.000000
R5_161 clk_6 clk_5 31.159999
R6_161 clk_6 clk_7 4.000000
R7_161 clk_7 clk 4.000000

C1_52 PNN130 0 0.004908PF
C2_52 PNN130_5 0 0.004929PF
C3_52 PNN130_4 0 0.000121PF
C4_52 PNN130_3 0 0.000189PF
C5_52 PNN130_2 0 0.000189PF
C6_52 iDFF_34_q_reg:D 0 0.000045PF
R1_52 iDFF_34_q_reg:D PNN130_2 4.000000
R2_52 PNN130_3 PNN130_2 1.976000
R3_52 PNN130_3 PNN130_4 4.000000
R4_52 PNN130_4 PNN130_5 4.000000
R5_52 PNN130 PNN130_5 45.143999

C1_219 U209:Z 0 0.000045PF
C2_219 n157_10 0 0.000035PF
C3_219 n157_9 0 0.000051PF
C4_219 n157_8 0 0.000727PF
C5_219 n157_7 0 0.000727PF
C6_219 n157_6 0 0.000043PF
C7_219 n157_5 0 0.000043PF
C8_219 n157_4 0 0.000242PF
C9_219 n157_3 0 0.000242PF
C10_219 n157_2 0 0.000121PF
C11_219 U207:A 0 0.000045PF
R1_219 U207:A n157_2 4.000000
R2_219 n157_2 n157_3 4.000000
R3_219 n157_3 n157_4 0.608000
R4_219 n157_4 n157_5 4.000000
R5_219 n157_6 n157_5 0.304000
R6_219 n157_6 n157_7 4.000000
R7_219 n157_7 n157_8 7.752000
R8_219 n157_8 n157_9 4.000000
R9_219 n157_9 n157_10 0.152000
R10_219 n157_10 U209:Z 4.000000

C1_137 oDFF_23_q_reg:Q 0 0.000045PF
C2_137 Qout_PNN746_8 0 0.000936PF
C3_137 Qout_PNN746_7 0 0.000936PF
C4_137 Qout_PNN746_6 0 0.000121PF
C5_137 Qout_PNN746_5 0 0.001895PF
C6_137 Qout_PNN746_4 0 0.001895PF
C7_137 Qout_PNN746_3 0 0.000044PF
C8_137 Qout_PNN746_2 0 0.000044PF
C9_137 Qout_PNN746 0 0.000042PF
R1_137 Qout_PNN746 Qout_PNN746_2 4.000000
R2_137 Qout_PNN746_3 Qout_PNN746_2 0.304000
R3_137 Qout_PNN746_3 Qout_PNN746_4 4.000000
R4_137 Qout_PNN746_5 Qout_PNN746_4 21.735999
R5_137 Qout_PNN746_5 Qout_PNN746_6 4.000000
R6_137 Qout_PNN746_6 Qout_PNN746_7 4.000000
R7_137 Qout_PNN746_8 Qout_PNN746_7 9.120000
R8_137 Qout_PNN746_8 oDFF_23_q_reg:Q 4.000000

C1_82 PNN97 0 0.000042PF
C2_82 PNN97_13 0 0.000121PF
C3_82 PNN97_12 0 0.000743PF
C4_82 PNN97_11 0 0.000743PF
C5_82 PNN97_10 0 0.000121PF
C6_82 PNN97_9 0 0.002402PF
C7_82 PNN97_8 0 0.002402PF
C8_82 PNN97_7 0 0.000121PF
C9_82 PNN97_6 0 0.000058PF
C10_82 PNN97_5 0 0.000058PF
C11_82 PNN97_4 0 0.000121PF
C12_82 PNN97_3 0 0.000466PF
C13_82 PNN97_2 0 0.000466PF
C14_82 iDFF_25_q_reg:D 0 0.000045PF
R1_82 iDFF_25_q_reg:D PNN97_2 4.000000
R2_82 PNN97_2 PNN97_3 5.776000
R3_82 PNN97_3 PNN97_4 4.000000
R4_82 PNN97_4 PNN97_5 4.000000
R5_82 PNN97_5 PNN97_6 0.608000
R6_82 PNN97_6 PNN97_7 4.000000
R7_82 PNN97_7 PNN97_8 4.000000
R8_82 PNN97_8 PNN97_9 27.055999
R9_82 PNN97_9 PNN97_10 4.000000
R10_82 PNN97_10 PNN97_11 4.000000
R11_82 PNN97_11 PNN97_12 7.600000
R12_82 PNN97_12 PNN97_13 4.000000
R13_82 PNN97_13 PNN97 4.000000

C1_65 PNN37 0 0.000042PF
C2_65 PNN37_15 0 0.000121PF
C3_65 PNN37_14 0 0.000814PF
C4_65 PNN37_13 0 0.000814PF
C5_65 PNN37_12 0 0.000121PF
C6_65 PNN37_11 0 0.002827PF
C7_65 PNN37_10 0 0.002827PF
C8_65 PNN37_9 0 0.000038PF
C9_65 PNN37_8 0 0.000055PF
C10_65 PNN37_7 0 0.001303PF
C11_65 PNN37_6 0 0.001303PF
C12_65 PNN37_5 0 0.000052PF
C13_65 PNN37_4 0 0.000036PF
C14_65 PNN37_3 0 0.000106PF
C15_65 PNN37_2 0 0.000106PF
C16_65 iDFF_10_q_reg:D 0 0.000045PF
R1_65 iDFF_10_q_reg:D PNN37_2 4.000000
R2_65 PNN37_3 PNN37_2 1.216000
R3_65 PNN37_3 PNN37_4 4.000000
R4_65 PNN37_5 PNN37_4 0.152000
R5_65 PNN37_5 PNN37_6 4.000000
R6_65 PNN37_7 PNN37_6 7.448000
R7_65 PNN37_7 PNN37_8 4.000000
R8_65 PNN37_8 PNN37_9 0.152000
R9_65 PNN37_9 PNN37_10 4.000000
R10_65 PNN37_11 PNN37_10 23.863999
R11_65 PNN37_11 PNN37_12 4.000000
R12_65 PNN37_12 PNN37_13 4.000000
R13_65 PNN37_14 PNN37_13 6.688000
R14_65 PNN37_14 PNN37_15 4.000000
R15_65 PNN37_15 PNN37 4.000000

C1_6 iDFF_29_q_reg:Q 0 0.000045PF
C2_6 INP_PNN113_16 0 0.000121PF
C3_6 INP_PNN113_13 0 0.000263PF
C4_6 INP_PNN113_11 0 0.000045PF
C5_6 INP_PNN113_9 0 0.000045PF
C6_6 INP_PNN113_7 0 0.001516PF
C7_6 INP_PNN113_5 0 0.001516PF
C8_6 INP_PNN113_2 0 0.000136PF
C9_6 INP_PNN113_4 0 0.000074PF
C10_6 INP_PNN113_6 0 0.002006PF
C11_6 INP_PNN113_8 0 0.002006PF
C12_6 INP_PNN113_10 0 0.000565PF
C13_6 INP_PNN113_12 0 0.000565PF
C14_6 clk_r_REG48_S2:D 0 0.000045PF
C15_6 U221:C 0 0.000045PF
C16_6 INP_PNN113_19 0 0.000041PF
C17_6 INP_PNN113_17 0 0.000041PF
C18_6 INP_PNN113_15 0 0.000263PF
C19_6 U199:C 0 0.000045PF
C20_6 INP_PNN113_1 0 0.000081PF
R1_6 INP_PNN113_1 INP_PNN113_2 0.608000
R2_6 INP_PNN113_1 U199:C 4.000000
R3_6 INP_PNN113_2 INP_PNN113_4 0.608000
R4_6 INP_PNN113_2 INP_PNN113_5 4.000000
R5_6 INP_PNN113_4 INP_PNN113_6 4.000000
R6_6 INP_PNN113_5 INP_PNN113_7 6.232000
R7_6 INP_PNN113_8 INP_PNN113_6 12.160000
R8_6 INP_PNN113_7 INP_PNN113_9 4.000000
R9_6 INP_PNN113_8 INP_PNN113_10 4.000000
R10_6 INP_PNN113_11 INP_PNN113_9 0.304000
R11_6 INP_PNN113_10 INP_PNN113_12 2.888000
R12_6 INP_PNN113_11 INP_PNN113_13 4.000000
R13_6 INP_PNN113_12 clk_r_REG48_S2:D 4.000000
R14_6 INP_PNN113_13 INP_PNN113_15 1.064000
R15_6 INP_PNN113_13 INP_PNN113_16 4.000000
R16_6 INP_PNN113_15 INP_PNN113_17 4.000000
R17_6 INP_PNN113_16 iDFF_29_q_reg:Q 4.000000
R18_6 INP_PNN113_19 INP_PNN113_17 0.304000
R19_6 INP_PNN113_19 U221:C 4.000000

C1_56 PNN134 0 0.003850PF
C2_56 PNN134_5 0 0.003871PF
C3_56 PNN134_4 0 0.000121PF
C4_56 PNN134_3 0 0.000170PF
C5_56 PNN134_2 0 0.000170PF
C6_56 iDFF_38_q_reg:D 0 0.000045PF
R1_56 iDFF_38_q_reg:D PNN134_2 4.000000
R2_56 PNN134_3 PNN134_2 1.672000
R3_56 PNN134_3 PNN134_4 4.000000
R4_56 PNN134_4 PNN134_5 4.000000
R5_56 PNN134 PNN134_5 47.119998

C1_133 oDFF_19_q_reg:Q 0 0.000045PF
C2_133 Qout_PNN742_8 0 0.002224PF
C3_133 Qout_PNN742_7 0 0.002224PF
C4_133 Qout_PNN742_6 0 0.000121PF
C5_133 Qout_PNN742_5 0 0.000576PF
C6_133 Qout_PNN742_4 0 0.000576PF
C7_133 Qout_PNN742_3 0 0.000044PF
C8_133 Qout_PNN742_2 0 0.000044PF
C9_133 Qout_PNN742 0 0.000042PF
R1_133 Qout_PNN742 Qout_PNN742_2 4.000000
R2_133 Qout_PNN742_3 Qout_PNN742_2 0.304000
R3_133 Qout_PNN742_3 Qout_PNN742_4 4.000000
R4_133 Qout_PNN742_5 Qout_PNN742_4 6.992000
R5_133 Qout_PNN742_5 Qout_PNN742_6 4.000000
R6_133 Qout_PNN742_6 Qout_PNN742_7 4.000000
R7_133 Qout_PNN742_8 Qout_PNN742_7 27.663999
R8_133 Qout_PNN742_8 oDFF_19_q_reg:Q 4.000000

C1_317 U286:B 0 0.000045PF
C2_317 n90_9 0 0.000033PF
C3_317 n90_8 0 0.000049PF
C4_317 n90_7 0 0.000121PF
C5_317 n90_6 0 0.000056PF
C6_317 n90_5 0 0.000056PF
C7_317 n90_4 0 0.000121PF
C8_317 n90_3 0 0.000071PF
C9_317 n90_2 0 0.000071PF
C10_317 U287:Z 0 0.000045PF
R1_317 U287:Z n90_2 4.000000
R2_317 n90_2 n90_3 0.608000
R3_317 n90_3 n90_4 4.000000
R4_317 n90_4 n90_5 4.000000
R5_317 n90_5 n90_6 0.760000
R6_317 n90_6 n90_7 4.000000
R7_317 n90_7 n90_8 4.000000
R8_317 n90_8 n90_9 0.152000
R9_317 n90_9 U286:B 4.000000

C1_1 FE_OFCC1_n168:Z 0 0.000046PF
C2_1 FE_OFCN1_n168_23 0 0.000068PF
C3_1 FE_OFCN1_n168_21 0 0.000568PF
C4_1 FE_OFCN1_n168_22 0 0.000530PF
C5_1 FE_OFCN1_n168_24 0 0.000826PF
C6_1 FE_OFCN1_n168_26 0 0.000826PF
C7_1 FE_OFCN1_n168_27 0 0.000063PF
C8_1 FE_OFCN1_n168_28 0 0.000063PF
C9_1 FE_OFCN1_n168_29 0 0.000617PF
C10_1 FE_OFCN1_n168_30 0 0.000617PF
C11_1 FE_OFCN1_n168_31 0 0.000060PF
C12_1 FE_OFCN1_n168_32 0 0.000060PF
C13_1 clk_r_REG25_S2:D 0 0.000045PF
C14_1 U168:B 0 0.000045PF
C15_1 FE_OFCN1_n168_15 0 0.000121PF
C16_1 FE_OFCN1_n168_13 0 0.000506PF
C17_1 FE_OFCN1_n168_14 0 0.000044PF
C18_1 FE_OFCN1_n168_16 0 0.000044PF
C19_1 FE_OFCN1_n168_18 0 0.000768PF
C20_1 FE_OFCN1_n168_19 0 0.000768PF
C21_1 FE_OFCN1_n168_20 0 0.000074PF
C22_1 U182:A 0 0.000045PF
C23_1 FE_OFCN1_n168_8 0 0.000767PF
C24_1 FE_OFCN1_n168_10 0 0.000506PF
C25_1 U166:A 0 0.000045PF
C26_1 FE_OFCN1_n168_9 0 0.000055PF
C27_1 FE_OFCN1_n168_7 0 0.000071PF
C28_1 FE_OFCN1_n168_4 0 0.000348PF
C29_1 FE_OFCN1_n168_2 0 0.000386PF
C30_1 FE_OFCN1_n168_5 0 0.000767PF
C31_1 U186:A 0 0.000045PF
C32_1 FE_OFCN1_n168_3 0 0.000121PF
C33_1 FE_OFCN1_n168_1 0 0.000057PF
R1_1 FE_OFCN1_n168_1 FE_OFCN1_n168_2 0.304000
R2_1 FE_OFCN1_n168_1 FE_OFCN1_n168_3 4.000000
R3_1 FE_OFCN1_n168_2 FE_OFCN1_n168_4 2.584000
R4_1 FE_OFCN1_n168_2 FE_OFCN1_n168_5 4.000000
R5_1 FE_OFCN1_n168_3 U186:A 4.000000
R6_1 FE_OFCN1_n168_4 FE_OFCN1_n168_7 4.000000
R7_1 FE_OFCN1_n168_5 FE_OFCN1_n168_8 3.952000
R8_1 FE_OFCN1_n168_7 FE_OFCN1_n168_9 0.152000
R9_1 FE_OFCN1_n168_8 FE_OFCN1_n168_10 4.000000
R10_1 FE_OFCN1_n168_8 U182:A 4.000000
R11_1 FE_OFCN1_n168_9 U166:A 4.000000
R12_1 FE_OFCN1_n168_10 FE_OFCN1_n168_13 3.648000
R13_1 FE_OFCN1_n168_13 FE_OFCN1_n168_14 4.000000
R14_1 FE_OFCN1_n168_13 FE_OFCN1_n168_15 4.000000
R15_1 FE_OFCN1_n168_16 FE_OFCN1_n168_14 0.304000
R16_1 FE_OFCN1_n168_15 U168:B 4.000000
R17_1 FE_OFCN1_n168_16 FE_OFCN1_n168_18 4.000000
R18_1 FE_OFCN1_n168_18 FE_OFCN1_n168_19 5.320000
R19_1 FE_OFCN1_n168_19 FE_OFCN1_n168_20 4.000000
R20_1 FE_OFCN1_n168_20 FE_OFCN1_n168_21 0.152000
R21_1 FE_OFCN1_n168_21 FE_OFCN1_n168_22 2.128000
R22_1 FE_OFCN1_n168_21 FE_OFCN1_n168_23 4.000000
R23_1 FE_OFCN1_n168_22 FE_OFCN1_n168_24 4.000000
R24_1 FE_OFCN1_n168_23 FE_OFCC1_n168:Z 0.456000
R25_1 FE_OFCN1_n168_24 FE_OFCN1_n168_26 3.496000
R26_1 FE_OFCN1_n168_26 FE_OFCN1_n168_27 4.000000
R27_1 FE_OFCN1_n168_27 FE_OFCN1_n168_28 0.608000
R28_1 FE_OFCN1_n168_28 FE_OFCN1_n168_29 4.000000
R29_1 FE_OFCN1_n168_29 FE_OFCN1_n168_30 6.536000
R30_1 FE_OFCN1_n168_30 FE_OFCN1_n168_31 4.000000
R31_1 FE_OFCN1_n168_32 FE_OFCN1_n168_31 0.304000
R32_1 FE_OFCN1_n168_32 clk_r_REG25_S2:D 4.000000

C1_199 U159:A 0 0.000045PF
C2_199 n137_4 0 0.000092PF
C3_199 n137_2 0 0.000970PF
C4_199 n137_5 0 0.000432PF
C5_199 n137_8 0 0.000432PF
C6_199 n137_10 0 0.000047PF
C7_199 n137_12 0 0.000047PF
C8_199 n137_14 0 0.000470PF
C9_199 n137_15 0 0.000504PF
C10_199 n137_16 0 0.001144PF
C11_199 n137_17 0 0.001110PF
C12_199 n137_18 0 0.000121PF
C13_199 U236:A 0 0.000095PF
C14_199 U254:Z 0 0.000045PF
C15_199 n137_11 0 0.000032PF
C16_199 n137_9 0 0.000049PF
C17_199 n137_6 0 0.000353PF
C18_199 n137_3 0 0.000353PF
C19_199 n137_1 0 0.000897PF
R1_199 n137_2 n137_1 10.488000
R2_199 n137_1 n137_3 4.000000
R3_199 n137_4 n137_2 1.368000
R4_199 n137_2 n137_5 4.000000
R5_199 n137_3 n137_6 0.912000
R6_199 n137_4 U159:A 4.000000
R7_199 n137_8 n137_5 2.584000
R8_199 n137_6 n137_9 4.000000
R9_199 n137_8 n137_10 4.000000
R10_199 n137_9 n137_11 0.152000
R11_199 n137_10 n137_12 0.304000
R12_199 n137_11 U254:Z 4.000000
R13_199 n137_12 n137_14 4.000000
R14_199 n137_15 n137_14 3.800000
R15_199 n137_16 n137_15 0.152000
R16_199 n137_17 n137_16 8.360000
R17_199 n137_17 n137_18 4.000000
R18_199 n137_18 U236:A 2.000000

C1_230 U187:A 0 0.000045PF
C2_230 n167_19 0 0.000121PF
C3_230 n167_17 0 0.000565PF
C4_230 n167_15 0 0.000565PF
C5_230 n167_12 0 0.000045PF
C6_230 n167_9 0 0.000258PF
C7_230 U183:C 0 0.000045PF
C8_230 U220:Z 0 0.000045PF
C9_230 n167_8 0 0.000121PF
C10_230 n167_4 0 0.003601PF
C11_230 n167_2 0 0.003687PF
C12_230 n167_5 0 0.000232PF
C13_230 clk_r_REG13_S2:D 0 0.000045PF
C14_230 n167_20 0 0.000055PF
C15_230 n167_18 0 0.000071PF
C16_230 n167_16 0 0.000475PF
C17_230 n167_14 0 0.000475PF
C18_230 n167_10 0 0.000045PF
C19_230 n167_7 0 0.000045PF
C20_230 U166:E 0 0.000045PF
C21_230 n167_3 0 0.000121PF
C22_230 n167_1 0 0.000104PF
R1_230 n167_1 n167_2 0.304000
R2_230 n167_1 n167_3 4.000000
R3_230 n167_2 n167_4 11.552000
R4_230 n167_2 n167_5 4.000000
R5_230 n167_3 U166:E 4.000000
R6_230 n167_4 n167_7 4.000000
R7_230 n167_4 n167_8 4.000000
R8_230 n167_9 n167_5 1.368000
R9_230 n167_10 n167_7 0.304000
R10_230 n167_8 U220:Z 4.000000
R11_230 n167_12 n167_9 0.304000
R12_230 n167_9 U183:C 4.000000
R13_230 n167_10 n167_14 4.000000
R14_230 n167_12 n167_15 4.000000
R15_230 n167_14 n167_16 2.736000
R16_230 n167_17 n167_15 2.584000
R17_230 n167_16 n167_18 4.000000
R18_230 n167_17 n167_19 4.000000
R19_230 n167_18 n167_20 0.152000
R20_230 n167_19 U187:A 4.000000
R21_230 n167_20 clk_r_REG13_S2:D 4.000000

C1_153 U233:A 0 0.000045PF
C2_153 c0_n31_13 0 0.000121PF
C3_153 c0_n31_9 0 0.001079PF
C4_153 c0_n31_5 0 0.001352PF
C5_153 c0_n31_2 0 0.000697PF
C6_153 c0_n31_4 0 0.000117PF
C7_153 c0_n31_7 0 0.000121PF
C8_153 c0_n31_11 0 0.000116PF
C9_153 c0_n31_15 0 0.000116PF
C10_153 clk_r_REG19_S2:D 0 0.000045PF
C11_153 U169:C 0 0.000045PF
C12_153 c0_n31_36 0 0.000121PF
C13_153 c0_n31_33 0 0.000121PF
C14_153 c0_n31_31 0 0.000064PF
C15_153 c0_n31_29 0 0.000064PF
C16_153 c0_n31_27 0 0.002952PF
C17_153 c0_n31_26 0 0.002517PF
C18_153 c0_n31_25 0 0.000213PF
C19_153 c0_n31_24 0 0.000213PF
C20_153 c0_n31_23 0 0.000326PF
C21_153 c0_n31_21 0 0.000326PF
C22_153 c0_n31_16 0 0.000125PF
C23_153 c0_n31_12 0 0.000110PF
C24_153 c0_n31_8 0 0.000291PF
C25_153 U188:A 0 0.000045PF
C26_153 c0_n31_32 0 0.000852PF
C27_153 c0_n31_30 0 0.000311PF
C28_153 c0_n31_28 0 0.000453PF
C29_153 U184:C 0 0.000045PF
C30_153 c0_n31_34 0 0.000559PF
C31_153 U173:Z 0 0.000045PF
C32_153 c0_n31_20 0 0.000034PF
C33_153 U245:A 0 0.000045PF
C34_153 c0_n31_14 0 0.000051PF
C35_153 c0_n31_10 0 0.000051PF
C36_153 c0_n31_6 0 0.000193PF
C37_153 c0_n31_3 0 0.000193PF
C38_153 c0_n31_1 0 0.000598PF
R1_153 c0_n31_2 c0_n31_1 7.296000
R2_153 c0_n31_1 c0_n31_3 4.000000
R3_153 c0_n31_4 c0_n31_2 1.216000
R4_153 c0_n31_2 c0_n31_5 4.000000
R5_153 c0_n31_3 c0_n31_6 2.128000
R6_153 c0_n31_4 c0_n31_7 4.000000
R7_153 c0_n31_8 c0_n31_5 3.192000
R8_153 c0_n31_5 c0_n31_9 4.712000
R9_153 c0_n31_6 c0_n31_10 4.000000
R10_153 c0_n31_7 c0_n31_11 4.000000
R11_153 c0_n31_8 c0_n31_12 4.000000
R12_153 c0_n31_9 c0_n31_13 4.000000
R13_153 c0_n31_10 c0_n31_14 0.304000
R14_153 c0_n31_15 c0_n31_11 1.216000
R15_153 c0_n31_12 c0_n31_16 1.064000
R16_153 c0_n31_13 U233:A 4.000000
R17_153 c0_n31_14 U245:A 4.000000
R18_153 c0_n31_15 clk_r_REG19_S2:D 4.000000
R19_153 c0_n31_16 c0_n31_20 0.152000
R20_153 c0_n31_16 c0_n31_21 4.000000
R21_153 c0_n31_20 U173:Z 4.000000
R22_153 c0_n31_23 c0_n31_21 1.368000
R23_153 c0_n31_23 c0_n31_24 4.000000
R24_153 c0_n31_24 c0_n31_25 0.912000
R25_153 c0_n31_25 c0_n31_26 4.000000
R26_153 c0_n31_27 c0_n31_26 10.640000
R27_153 c0_n31_28 c0_n31_27 1.672000
R28_153 c0_n31_27 c0_n31_29 4.000000
R29_153 c0_n31_28 c0_n31_30 4.000000
R30_153 c0_n31_31 c0_n31_29 0.456000
R31_153 c0_n31_30 c0_n31_32 3.648000
R32_153 c0_n31_31 c0_n31_33 4.000000
R33_153 c0_n31_32 c0_n31_34 3.952000
R34_153 c0_n31_32 U188:A 4.000000
R35_153 c0_n31_33 c0_n31_36 4.000000
R36_153 c0_n31_34 U184:C 4.000000
R37_153 c0_n31_36 U169:C 4.000000

C1_326 U305:B 0 0.000045PF
C2_326 n99_16 0 0.000121PF
C3_326 n99_13 0 0.001066PF
C4_326 n99_15 0 0.000138PF
C5_326 n99_18 0 0.000138PF
C6_326 n99_21 0 0.000506PF
C7_326 n99_22 0 0.000506PF
C8_326 n99_23 0 0.000272PF
C9_326 n99_24 0 0.000272PF
C10_326 U303:B 0 0.000045PF
C11_326 U301:B 0 0.000045PF
C12_326 n99_8 0 0.000121PF
C13_326 n99_4 0 0.001156PF
C14_326 n99_7 0 0.000156PF
C15_326 n99_10 0 0.001101PF
C16_326 U211:Z 0 0.000045PF
C17_326 n99_17 0 0.000076PF
C18_326 n99_14 0 0.000076PF
C19_326 n99_12 0 0.000121PF
C20_326 n99_9 0 0.000595PF
C21_326 n99_5 0 0.000595PF
C22_326 n99_2 0 0.001276PF
C23_326 U307:B 0 0.000045PF
C24_326 n99_3 0 0.000121PF
C25_326 n99_1 0 0.000241PF
R1_326 n99_1 n99_2 3.192000
R2_326 n99_1 n99_3 4.000000
R3_326 n99_2 n99_4 5.168000
R4_326 n99_2 n99_5 4.000000
R5_326 n99_3 U307:B 4.000000
R6_326 n99_4 n99_7 0.456000
R7_326 n99_4 n99_8 4.000000
R8_326 n99_5 n99_9 7.752000
R9_326 n99_10 n99_7 0.152000
R10_326 n99_8 U301:B 4.000000
R11_326 n99_9 n99_12 4.000000
R12_326 n99_10 n99_13 6.688000
R13_326 n99_12 n99_14 4.000000
R14_326 n99_13 n99_15 4.000000
R15_326 n99_13 n99_16 4.000000
R16_326 n99_14 n99_17 1.064000
R17_326 n99_18 n99_15 0.608000
R18_326 n99_16 U305:B 4.000000
R19_326 n99_17 U211:Z 4.000000
R20_326 n99_18 n99_21 4.000000
R21_326 n99_21 n99_22 4.408000
R22_326 n99_22 n99_23 4.000000
R23_326 n99_24 n99_23 2.128000
R24_326 n99_24 U303:B 4.000000

C1_79 PNN89 0 0.000042PF
C2_79 PNN89_7 0 0.000121PF
C3_79 PNN89_6 0 0.000668PF
C4_79 PNN89_5 0 0.000668PF
C5_79 PNN89_4 0 0.000121PF
C6_79 PNN89_3 0 0.002147PF
C7_79 PNN89_2 0 0.002147PF
C8_79 iDFF_23_q_reg:D 0 0.000045PF
R1_79 iDFF_23_q_reg:D PNN89_2 4.000000
R2_79 PNN89_2 PNN89_3 25.383999
R3_79 PNN89_3 PNN89_4 4.000000
R4_79 PNN89_4 PNN89_5 4.000000
R5_79 PNN89_5 PNN89_6 7.752000
R6_79 PNN89_6 PNN89_7 4.000000
R7_79 PNN89_7 PNN89 4.000000

C1_73 PNN65 0 0.004051PF
C2_73 PNN65_8 0 0.004072PF
C3_73 PNN65_7 0 0.000121PF
C4_73 PNN65_6 0 0.000283PF
C5_73 PNN65_5 0 0.000283PF
C6_73 PNN65_4 0 0.000121PF
C7_73 PNN65_3 0 0.000180PF
C8_73 PNN65_2 0 0.000180PF
C9_73 iDFF_17_q_reg:D 0 0.000045PF
R1_73 iDFF_17_q_reg:D PNN65_2 4.000000
R2_73 PNN65_2 PNN65_3 1.976000
R3_73 PNN65_3 PNN65_4 4.000000
R4_73 PNN65_4 PNN65_5 4.000000
R5_73 PNN65_5 PNN65_6 2.280000
R6_73 PNN65_6 PNN65_7 4.000000
R7_73 PNN65_7 PNN65_8 4.000000
R8_73 PNN65_8 PNN65 36.783999

C1_75 PNN73 0 0.002357PF
C2_75 PNN73_8 0 0.002378PF
C3_75 PNN73_7 0 0.000049PF
C4_75 PNN73_6 0 0.000033PF
C5_75 PNN73_5 0 0.001446PF
C6_75 PNN73_4 0 0.001481PF
C7_75 PNN73_3 0 0.000167PF
C8_75 PNN73_2 0 0.000133PF
C9_75 iDFF_19_q_reg:D 0 0.000045PF
R1_75 iDFF_19_q_reg:D PNN73_2 4.000000
R2_75 PNN73_2 PNN73_3 1.368000
R3_75 PNN73_3 PNN73_4 0.152000
R4_75 PNN73_4 PNN73_5 7.448000
R5_75 PNN73_5 PNN73_6 4.000000
R6_75 PNN73_7 PNN73_6 0.152000
R7_75 PNN73_7 PNN73_8 4.000000
R8_75 PNN73_8 PNN73 29.943999

C1_76 PNN77 0 0.000042PF
C2_76 PNN77_7 0 0.000121PF
C3_76 PNN77_6 0 0.000634PF
C4_76 PNN77_5 0 0.000634PF
C5_76 PNN77_4 0 0.000121PF
C6_76 PNN77_3 0 0.002098PF
C7_76 PNN77_2 0 0.002098PF
C8_76 iDFF_20_q_reg:D 0 0.000045PF
R1_76 iDFF_20_q_reg:D PNN77_2 4.000000
R2_76 PNN77_2 PNN77_3 25.383999
R3_76 PNN77_3 PNN77_4 4.000000
R4_76 PNN77_4 PNN77_5 4.000000
R5_76 PNN77_5 PNN77_6 7.752000
R6_76 PNN77_6 PNN77_7 4.000000
R7_76 PNN77_7 PNN77 4.000000

C1_30 clk_r_REG34_S2:D 0 0.000045PF
C2_30 INP_PNN57_14 0 0.000271PF
C3_30 INP_PNN57_13 0 0.000387PF
C4_30 INP_PNN57_12 0 0.000387PF
C5_30 INP_PNN57_10 0 0.000045PF
C6_30 INP_PNN57_7 0 0.000045PF
C7_30 INP_PNN57_4 0 0.000093PF
C8_30 INP_PNN57_2 0 0.000950PF
C9_30 INP_PNN57_5 0 0.000218PF
C10_30 INP_PNN57_8 0 0.000265PF
C11_30 U198:B 0 0.000095PF
C12_30 iDFF_15_q_reg:Q 0 0.000045PF
C13_30 INP_PNN57_20 0 0.000079PF
C14_30 INP_PNN57_19 0 0.000079PF
C15_30 INP_PNN57_18 0 0.000192PF
C16_30 INP_PNN57_17 0 0.000192PF
C17_30 INP_PNN57_15 0 0.000255PF
C18_30 U253:B 0 0.000045PF
C19_30 INP_PNN57_6 0 0.000058PF
C20_30 INP_PNN57_3 0 0.000058PF
C21_30 INP_PNN57_1 0 0.000875PF
R1_30 INP_PNN57_1 INP_PNN57_2 4.104000
R2_30 INP_PNN57_1 INP_PNN57_3 4.000000
R3_30 INP_PNN57_2 INP_PNN57_4 0.912000
R4_30 INP_PNN57_2 INP_PNN57_5 4.000000
R5_30 INP_PNN57_6 INP_PNN57_3 0.608000
R6_30 INP_PNN57_4 INP_PNN57_7 4.000000
R7_30 INP_PNN57_5 INP_PNN57_8 3.344000
R8_30 INP_PNN57_6 U253:B 4.000000
R9_30 INP_PNN57_10 INP_PNN57_7 0.304000
R10_30 INP_PNN57_8 U198:B 2.000000
R11_30 INP_PNN57_10 INP_PNN57_12 4.000000
R12_30 INP_PNN57_12 INP_PNN57_13 2.888000
R13_30 INP_PNN57_13 INP_PNN57_14 4.000000
R14_30 INP_PNN57_15 INP_PNN57_14 1.064000
R15_30 INP_PNN57_14 clk_r_REG34_S2:D 4.000000
R16_30 INP_PNN57_15 INP_PNN57_17 4.000000
R17_30 INP_PNN57_17 INP_PNN57_18 1.976000
R18_30 INP_PNN57_18 INP_PNN57_19 4.000000
R19_30 INP_PNN57_20 INP_PNN57_19 0.760000
R20_30 INP_PNN57_20 iDFF_15_q_reg:Q 4.000000

C1_71 PNN57 0 0.002298PF
C2_71 PNN57_5 0 0.002319PF
C3_71 PNN57_4 0 0.000121PF
C4_71 PNN57_3 0 0.000575PF
C5_71 PNN57_2 0 0.000575PF
C6_71 iDFF_15_q_reg:D 0 0.000045PF
R1_71 iDFF_15_q_reg:D PNN57_2 4.000000
R2_71 PNN57_3 PNN57_2 2.736000
R3_71 PNN57_3 PNN57_4 4.000000
R4_71 PNN57_4 PNN57_5 4.000000
R5_71 PNN57 PNN57_5 30.247999

C1_315 U202:Z 0 0.000251PF
C2_315 n89_40 0 0.000274PF
C3_315 n89_39 0 0.000564PF
C4_315 n89_38 0 0.000564PF
C5_315 n89_37 0 0.000904PF
C6_315 n89_36 0 0.000904PF
C7_315 n89_35 0 0.000110PF
C8_315 n89_34 0 0.000110PF
C9_315 n89_33 0 0.000121PF
C10_315 n89_32 0 0.000121PF
C11_315 n89_31 0 0.000069PF
C12_315 n89_30 0 0.000069PF
C13_315 n89_29 0 0.002555PF
C14_315 n89_27 0 0.002555PF
C15_315 n89_25 0 0.000406PF
C16_315 n89_26 0 0.000377PF
C17_315 U287:B 0 0.000045PF
C18_315 U289:B 0 0.000045PF
C19_315 n89_19 0 0.000136PF
C20_315 n89_15 0 0.000136PF
C21_315 n89_11 0 0.000121PF
C22_315 n89_7 0 0.000079PF
C23_315 n89_4 0 0.000127PF
C24_315 n89_8 0 0.001414PF
C25_315 n89_12 0 0.001414PF
C26_315 n89_16 0 0.000056PF
C27_315 n89_20 0 0.000056PF
C28_315 n89_22 0 0.000062PF
C29_315 n89_23 0 0.000062PF
C30_315 n89_24 0 0.000047PF
C31_315 U291:B 0 0.000045PF
C32_315 n89_13 0 0.000121PF
C33_315 n89_9 0 0.000049PF
C34_315 n89_5 0 0.000049PF
C35_315 n89_2 0 0.000127PF
C36_315 U285:B 0 0.000045PF
C37_315 n89_14 0 0.000328PF
C38_315 n89_10 0 0.000328PF
C39_315 n89_6 0 0.000051PF
C40_315 n89_3 0 0.000051PF
C41_315 n89_1 0 0.000079PF
R1_315 n89_2 n89_1 0.760000
R2_315 n89_1 n89_3 4.000000
R3_315 n89_4 n89_2 0.608000
R4_315 n89_2 n89_5 4.000000
R5_315 n89_3 n89_6 0.304000
R6_315 n89_7 n89_4 0.760000
R7_315 n89_4 n89_8 4.000000
R8_315 n89_9 n89_5 0.304000
R9_315 n89_6 n89_10 4.000000
R10_315 n89_7 n89_11 4.000000
R11_315 n89_12 n89_8 9.120000
R12_315 n89_9 n89_13 4.000000
R13_315 n89_10 n89_14 4.256000
R14_315 n89_11 n89_15 4.000000
R15_315 n89_12 n89_16 4.000000
R16_315 n89_13 U291:B 4.000000
R17_315 n89_14 U285:B 4.000000
R18_315 n89_19 n89_15 2.432000
R19_315 n89_16 n89_20 0.456000
R20_315 n89_19 U289:B 4.000000
R21_315 n89_20 n89_22 4.000000
R22_315 n89_23 n89_22 0.456000
R23_315 n89_23 n89_24 4.000000
R24_315 n89_24 n89_25 0.304000
R25_315 n89_25 n89_26 3.648000
R26_315 n89_25 n89_27 4.000000
R27_315 n89_26 U287:B 4.000000
R28_315 n89_29 n89_27 9.728000
R29_315 n89_29 n89_30 4.000000
R30_315 n89_31 n89_30 0.456000
R31_315 n89_31 n89_32 4.000000
R32_315 n89_33 n89_32 0.456000
R33_315 n89_33 n89_34 4.000000
R34_315 n89_35 n89_34 0.304000
R35_315 n89_35 n89_36 4.000000
R36_315 n89_37 n89_36 5.320000
R37_315 n89_37 n89_38 4.000000
R38_315 n89_39 n89_38 5.320000
R39_315 n89_39 n89_40 4.000000
R40_315 U202:Z n89_40 2.432000

C1_125 oDFF_11_q_reg:Q 0 0.000045PF
C2_125 Qout_PNN734_9 0 0.003502PF
C3_125 Qout_PNN734_8 0 0.003502PF
C4_125 Qout_PNN734_7 0 0.000136PF
C5_125 Qout_PNN734_6 0 0.000136PF
C6_125 Qout_PNN734_5 0 0.000045PF
C7_125 Qout_PNN734_4 0 0.000045PF
C8_125 Qout_PNN734_3 0 0.000079PF
C9_125 Qout_PNN734_2 0 0.000079PF
C10_125 Qout_PNN734 0 0.000042PF
R1_125 Qout_PNN734 Qout_PNN734_2 4.000000
R2_125 Qout_PNN734_2 Qout_PNN734_3 0.760000
R3_125 Qout_PNN734_3 Qout_PNN734_4 4.000000
R4_125 Qout_PNN734_4 Qout_PNN734_5 0.304000
R5_125 Qout_PNN734_5 Qout_PNN734_6 4.000000
R6_125 Qout_PNN734_6 Qout_PNN734_7 1.520000
R7_125 Qout_PNN734_7 Qout_PNN734_8 4.000000
R8_125 Qout_PNN734_8 Qout_PNN734_9 30.399999
R9_125 Qout_PNN734_9 oDFF_11_q_reg:Q 4.000000

C1_162 iDFF_24_q_reg:CP 0 0.000045PF
C2_162 clk__L1_N0_64 0 0.000121PF
C3_162 clk__L1_N0_56 0 0.000442PF
C4_162 clk__L1_N0_48 0 0.000794PF
C5_162 clk__L1_N0_57 0 0.000194PF
C6_162 clk__L1_N0_65 0 0.000194PF
C7_162 clk__L1_N0_74 0 0.000121PF
C8_162 clk__L1_N0_82 0 0.000121PF
C9_162 oDFF_20_q_reg:CP 0 0.000045PF
C10_162 iDFF_20_q_reg:CP 0 0.000045PF
C11_162 clk__L1_N0_49 0 0.000121PF
C12_162 clk__L1_N0_39 0 0.000531PF
C13_162 iDFF_23_q_reg:CP 0 0.000045PF
C14_162 clk__L1_N0_40 0 0.000121PF
C15_162 clk__L1_N0_31 0 0.000245PF
C16_162 clk_r_REG42_S2:CP 0 0.000045PF
C17_162 clk__L1_N0_32 0 0.000121PF
C18_162 clk__L1_N0_25 0 0.000085PF
C19_162 oDFF_19_q_reg:CP 0 0.000045PF
C20_162 clk__L1_N0_17 0 0.000121PF
C21_162 clk__L1_N0_11 0 0.000481PF
C22_162 clk__L1_N0_7 0 0.000700PF
C23_162 clk__L1_N0_4 0 0.000257PF
C24_162 clk__L1_N0_2 0 0.000329PF
C25_162 clk__L1_N0_5 0 0.000281PF
C26_162 clk__L1_N0_8 0 0.000281PF
C27_162 clk__L1_N0_12 0 0.000129PF
C28_162 clk__L1_N0_18 0 0.000129PF
C29_162 clk_r_REG38_S2:CP 0 0.000045PF
C30_162 clk__L1_N0_47 0 0.000121PF
C31_162 clk__L1_N0_38 0 0.000121PF
C32_162 clk__L1_N0_30 0 0.000260PF
C33_162 clk__L1_N0_23 0 0.000260PF
C34_162 clk__L1_N0_16 0 0.000700PF
C35_162 clk_r_REG39_S2:CP 0 0.000045PF
C36_162 clk__L1_N0_29 0 0.000121PF
C37_162 clk__L1_N0_22 0 0.001060PF
C38_162 clk_r_REG43_S2:CP 0 0.000045PF
C39_162 clk__L1_N0_36 0 0.000121PF
C40_162 clk__L1_N0_28 0 0.000744PF
C41_162 oDFF_24_q_reg:CP 0 0.000045PF
C42_162 clk__L1_N0_72 0 0.000121PF
C43_162 clk__L1_N0_63 0 0.000095PF
C44_162 clk__L1_N0_54 0 0.000095PF
C45_162 clk__L1_N0_45 0 0.000194PF
C46_162 clk__L1_N0_35 0 0.000194PF
C47_162 iDFF_21_q_reg:CP 0 0.000045PF
C48_162 clk__L1_N0_102 0 0.000121PF
C49_162 clk__L1_N0_95 0 0.000180PF
C50_162 clk__L1_N0_88 0 0.000180PF
C51_162 clk__L1_N0_80 0 0.000148PF
C52_162 clk__L1_N0_71 0 0.000148PF
C53_162 iDFF_28_q_reg:CP 0 0.000045PF
C54_162 clk__L1_N0_15 0 0.000121PF
C55_162 clk__L1_N0_10 0 0.000638PF
C56_162 iDFF_32_q_reg:CP 0 0.000045PF
C57_162 clk__L1_N0_34 0 0.000121PF
C58_162 clk__L1_N0_27 0 0.000301PF
C59_162 clk__L1_N0_20 0 0.000109PF
C60_162 clk__L1_N0_14 0 0.000109PF
C61_162 iDFF_31_q_reg:CP 0 0.000045PF
C62_162 clk__L1_N0_43 0 0.000121PF
C63_162 clk__L1_N0_33 0 0.000310PF
C64_162 oDFF_28_q_reg:CP 0 0.000045PF
C65_162 clk__L1_N0_52 0 0.000121PF
C66_162 clk__L1_N0_42 0 0.000365PF
C67_162 clk_r_REG51_S2:CP 0 0.000045PF
C68_162 clk__L1_N0_61 0 0.000121PF
C69_162 clk__L1_N0_51 0 0.000672PF
C70_162 clk_r_REG50_S2:CP 0 0.000045PF
C71_162 clk__L1_N0_94 0 0.000121PF
C72_162 clk__L1_N0_87 0 0.000050PF
C73_162 clk__L1_N0_79 0 0.000050PF
C74_162 clk__L1_N0_69 0 0.000325PF
C75_162 clk__L1_N0_60 0 0.000149PF
C76_162 oDFF_27_q_reg:CP 0 0.000045PF
C77_162 clk__L1_N0_93 0 0.000121PF
C78_162 clk__L1_N0_86 0 0.000266PF
C79_162 clk__L1_N0_78 0 0.000317PF
C80_162 clk_r_REG44_S2:CP 0 0.000045PF
C81_162 clk__L1_N0_99 0 0.000121PF
C82_162 clk__L1_N0_92 0 0.000312PF
C83_162 iDFF_27_q_reg:CP 0 0.000045PF
C84_162 clk__L1_N0_121 0 0.000121PF
C85_162 clk__L1_N0_115 0 0.000125PF
C86_162 clk__L1_N0_111 0 0.000143PF
C87_162 clk__L1_N0_106 0 0.000153PF
C88_162 clk__L1_N0_98 0 0.000153PF
C89_162 clk_r_REG16_S2:CP 0 0.000045PF
C90_162 clk__L1_N0_158 0 0.000121PF
C91_162 clk__L1_N0_148 0 0.000439PF
C92_162 clk__L1_N0_138 0 0.000060PF
C93_162 clk__L1_N0_128 0 0.000183PF
C94_162 clk__L1_N0_120 0 0.000183PF
C95_162 iDFF_29_q_reg:CP 0 0.000045PF
C96_162 clk__L1_N0_203 0 0.000121PF
C97_162 clk__L1_N0_197 0 0.000121PF
C98_162 clk__L1_N0_190 0 0.000097PF
C99_162 clk__L1_N0_183 0 0.000097PF
C100_162 clk__L1_N0_175 0 0.000172PF
C101_162 clk__L1_N0_166 0 0.000109PF
C102_162 clk__L1_N0_157 0 0.000433PF
C103_162 iDFF_25_q_reg:CP 0 0.000045PF
C104_162 clk__L1_N0_189 0 0.000121PF
C105_162 clk__L1_N0_182 0 0.000600PF
C106_162 iDFF_17_q_reg:CP 0 0.000045PF
C107_162 clk__L1_N0_195 0 0.000121PF
C108_162 clk__L1_N0_188 0 0.000503PF
C109_162 iDFF_19_q_reg:CP 0 0.000045PF
C110_162 clk__L1_N0_215 0 0.000121PF
C111_162 clk__L1_N0_208 0 0.000430PF
C112_162 clk__L1_N0_201 0 0.000223PF
C113_162 clk__L1_N0_194 0 0.000223PF
C114_162 clk_r_REG25_S2:CP 0 0.000045PF
C115_162 clk__L1_N0_231 0 0.000055PF
C116_162 clk__L1_N0_222 0 0.000071PF
C117_162 clk__L1_N0_214 0 0.000575PF
C118_162 clk_r_REG36_S2:CP 0 0.000045PF
C119_162 clk__L1_N0_250 0 0.000121PF
C120_162 clk__L1_N0_244 0 0.000078PF
C121_162 clk__L1_N0_238 0 0.000078PF
C122_162 clk__L1_N0_230 0 0.000201PF
C123_162 clk__L1_N0_221 0 0.000201PF
C124_162 clk_r_REG40_S2:CP 0 0.000045PF
C125_162 clk__L1_N0_229 0 0.000121PF
C126_162 clk__L1_N0_220 0 0.000422PF
C127_162 oDFF_17_q_reg:CP 0 0.000045PF
C128_162 clk__L1_N0_236 0 0.000121PF
C129_162 clk__L1_N0_228 0 0.000344PF
C130_162 oDFF_21_q_reg:CP 0 0.000045PF
C131_162 clk__L1_N0_271 0 0.000121PF
C132_162 clk__L1_N0_264 0 0.000117PF
C133_162 clk__L1_N0_257 0 0.000117PF
C134_162 clk__L1_N0_249 0 0.000321PF
C135_162 clk__L1_N0_242 0 0.000321PF
C136_162 clk__L1_N0_235 0 0.000103PF
C137_162 clk_r_REG46_S2:CP 0 0.000045PF
C138_162 clk__L1_N0_119 0 0.000121PF
C139_162 clk__L1_N0_114 0 0.000036PF
C140_162 clk_r_REG24_S2:CP 0 0.000045PF
C141_162 clk__L1_N0_105 0 0.000121PF
C142_162 clk__L1_N0_97 0 0.000428PF
C143_162 clk__L1_N0_91 0 0.000412PF
C144_162 clk__L1_N0_85 0 0.000141PF
C145_162 clk_r_REG15_S2:CP 0 0.000045PF
C146_162 clk__L1_N0_126 0 0.000121PF
C147_162 clk__L1_N0_118 0 0.000039PF
C148_162 clk__L1_N0_113 0 0.000291PF
C149_162 clk__L1_N0_109 0 0.000249PF
C150_162 clk__L1_N0_104 0 0.000206PF
C151_162 clk_r_REG12_S2:CP 0 0.000045PF
C152_162 clk__L1_N0_136 0 0.000036PF
C153_162 clk__L1_N0_125 0 0.000052PF
C154_162 clk__L1_N0_117 0 0.000605PF
C155_162 iDFF_26_q_reg:CP 0 0.000045PF
C156_162 clk__L1_N0_135 0 0.000121PF
C157_162 clk__L1_N0_124 0 0.000414PF
C158_162 clk_r_REG49_S2:CP 0 0.000045PF
C159_162 clk__L1_N0_174 0 0.000121PF
C160_162 clk__L1_N0_165 0 0.000217PF
C161_162 clk__L1_N0_156 0 0.000217PF
C162_162 clk__L1_N0_145 0 0.000102PF
C163_162 clk__L1_N0_134 0 0.000285PF
C164_162 clk_r_REG48_S2:CP 0 0.000045PF
C165_162 clk__L1_N0_173 0 0.000121PF
C166_162 clk__L1_N0_164 0 0.000188PF
C167_162 clk__L1_N0_155 0 0.000188PF
C168_162 clk__L1_N0_144 0 0.000201PF
C169_162 oDFF_26_q_reg:CP 0 0.000045PF
C170_162 clk__L1_N0_143 0 0.000121PF
C171_162 clk__L1_N0_133 0 0.000232PF
C172_162 oDFF_29_q_reg:CP 0 0.000045PF
C173_162 clk__L1_N0_179 0 0.000121PF
C174_162 clk__L1_N0_172 0 0.000121PF
C175_162 clk__L1_N0_163 0 0.000328PF
C176_162 clk__L1_N0_153 0 0.000328PF
C177_162 clk__L1_N0_142 0 0.000206PF
C178_162 iDFF_30_q_reg:CP 0 0.000045PF
C179_162 clk__L1_N0_186 0 0.000121PF
C180_162 clk__L1_N0_178 0 0.000121PF
C181_162 clk__L1_N0_171 0 0.000153PF
C182_162 clk__L1_N0_162 0 0.000153PF
C183_162 clk__L1_N0_152 0 0.000056PF
C184_162 clk_r_REG45_S2:CP 0 0.000045PF
C185_162 clk__L1_N0_141 0 0.000061PF
C186_162 clk__L1_N0_132 0 0.000061PF
C187_162 clk__L1_N0_123 0 0.000121PF
C188_162 clk__L1_N0_116 0 0.000324PF
C189_162 clk__L1_N0_112 0 0.000160PF
C190_162 clk_r_REG27_S2:CP 0 0.000045PF
C191_162 clk__L1_N0_150 0 0.000121PF
C192_162 clk__L1_N0_140 0 0.000039PF
C193_162 clk__L1_N0_131 0 0.000055PF
C194_162 clk__L1_N0_122 0 0.000346PF
C195_162 clk_r_REG14_S2:CP 0 0.000045PF
C196_162 clk__L1_N0_160 0 0.000121PF
C197_162 clk__L1_N0_149 0 0.000808PF
C198_162 clk__L1_N0_139 0 0.000248PF
C199_162 clk__L1_N0_130 0 0.000148PF
C200_162 oDFF_30_q_reg:CP 0 0.000045PF
C201_162 clk__L1_N0_169 0 0.000121PF
C202_162 clk__L1_N0_159 0 0.000596PF
C203_162 clk_r_REG11_S2:CP 0 0.000045PF
C204_162 clk__L1_N0_200 0 0.000121PF
C205_162 clk__L1_N0_192 0 0.000121PF
C206_162 clk__L1_N0_185 0 0.000121PF
C207_162 clk__L1_N0_176 0 0.000497PF
C208_162 clk__L1_N0_168 0 0.000194PF
C209_162 clk_r_REG8_S2:CP 0 0.000045PF
C210_162 clk__L1_N0_227 0 0.000121PF
C211_162 clk__L1_N0_219 0 0.000195PF
C212_162 clk__L1_N0_213 0 0.000148PF
C213_162 clk__L1_N0_206 0 0.000148PF
C214_162 clk__L1_N0_199 0 0.000289PF
C215_162 clk__L1_N0_191 0 0.000196PF
C216_162 clk__L1_N0_184 0 0.000321PF
C217_162 oDFF_4_q_reg:CP 0 0.000045PF
C218_162 clk__L1_N0_256 0 0.000121PF
C219_162 clk__L1_N0_248 0 0.000121PF
C220_162 clk__L1_N0_241 0 0.000324PF
C221_162 clk__L1_N0_233 0 0.000183PF
C222_162 clk__L1_N0_226 0 0.000132PF
C223_162 clk_r_REG1_S2:CP 0 0.000045PF
C224_162 clk__L1_N0_270 0 0.000121PF
C225_162 clk__L1_N0_262 0 0.000374PF
C226_162 clk__L1_N0_255 0 0.000244PF
C227_162 clk__L1_N0_247 0 0.000331PF
C228_162 iDFF_1_q_reg:CP 0 0.000045PF
C229_162 clk__L1_N0_277 0 0.000121PF
C230_162 clk__L1_N0_269 0 0.000148PF
C231_162 iDFF_8_q_reg:CP 0 0.000045PF
C232_162 clk__L1_N0_285 0 0.000055PF
C233_162 clk__L1_N0_276 0 0.000071PF
C234_162 clk__L1_N0_268 0 0.000079PF
C235_162 clk__L1_N0_261 0 0.000094PF
C236_162 clk__L1_N0_254 0 0.000189PF
C237_162 oDFF_1_q_reg:CP 0 0.000045PF
C238_162 clk__L1_N0_275 0 0.000121PF
C239_162 clk__L1_N0_267 0 0.000071PF
C240_162 clk_r_REG7_S2:CP 0 0.000045PF
C241_162 clk__L1_N0_307 0 0.000121PF
C242_162 clk__L1_N0_301 0 0.000083PF
C243_162 clk__L1_N0_296 0 0.000083PF
C244_162 clk__L1_N0_290 0 0.000324PF
C245_162 clk__L1_N0_283 0 0.000160PF
C246_162 clk__L1_N0_274 0 0.000202PF
C247_162 oDFF_8_q_reg:CP 0 0.000045PF
C248_162 clk__L1_N0_306 0 0.000121PF
C249_162 clk__L1_N0_300 0 0.000220PF
C250_162 clk__L1_N0_295 0 0.000183PF
C251_162 clk_r_REG2_S2:CP 0 0.000045PF
C252_162 clk__L1_N0_327 0 0.000033PF
C253_162 clk__L1_N0_321 0 0.000049PF
C254_162 clk__L1_N0_317 0 0.000188PF
C255_162 clk__L1_N0_315 0 0.000147PF
C256_162 clk__L1_N0_310 0 0.000147PF
C257_162 clk__L1_N0_305 0 0.000203PF
C258_162 oDFF_5_q_reg:CP 0 0.000045PF
C259_162 clk__L1_N0_326 0 0.000121PF
C260_162 clk__L1_N0_320 0 0.000267PF
C261_162 iDFF_5_q_reg:CP 0 0.000045PF
C262_162 clk__L1_N0_355 0 0.000121PF
C263_162 clk__L1_N0_347 0 0.000121PF
C264_162 clk__L1_N0_340 0 0.000247PF
C265_162 clk__L1_N0_332 0 0.000090PF
C266_162 clk__L1_N0_325 0 0.000277PF
C267_162 clk_r_REG0_S2:CP 0 0.000045PF
C268_162 clk__L1_N0_377 0 0.000121PF
C269_162 clk__L1_N0_364 0 0.000157PF
C270_162 clk__L1_N0_354 0 0.000045PF
C271_162 clk__L1_N0_346 0 0.000176PF
C272_162 oDFF_9_q_reg:CP 0 0.000045PF
C273_162 clk__L1_N0_419 0 0.000121PF
C274_162 clk__L1_N0_408 0 0.000121PF
C275_162 clk__L1_N0_397 0 0.000141PF
C276_162 clk__L1_N0_387 0 0.000141PF
C277_162 clk__L1_N0_376 0 0.000131PF
C278_162 oDFF_13_q_reg:CP 0 0.000045PF
C279_162 clk__L1_N0_345 0 0.000055PF
C280_162 clk__L1_N0_339 0 0.000071PF
C281_162 clk__L1_N0_331 0 0.000396PF
C282_162 iDFF_13_q_reg:CP 0 0.000045PF
C283_162 clk__L1_N0_375 0 0.000121PF
C284_162 clk__L1_N0_363 0 0.000121PF
C285_162 clk__L1_N0_352 0 0.000312PF
C286_162 clk__L1_N0_344 0 0.000137PF
C287_162 clk__L1_N0_338 0 0.000303PF
C288_162 clk_r_REG23_S2:CP 0 0.000045PF
C289_162 clk__L1_N0_385 0 0.000121PF
C290_162 clk__L1_N0_374 0 0.000121PF
C291_162 clk__L1_N0_362 0 0.000315PF
C292_162 clk_r_REG26_S2:CP 0 0.000045PF
C293_162 clk__L1_N0_407 0 0.000121PF
C294_162 clk__L1_N0_395 0 0.000402PF
C295_162 clk__L1_N0_384 0 0.000310PF
C296_162 clk__L1_N0_373 0 0.000139PF
C297_162 iDFF_9_q_reg:CP 0 0.000045PF
C298_162 clk__L1_N0_417 0 0.000121PF
C299_162 clk__L1_N0_406 0 0.000417PF
C300_162 iDFF_12_q_reg:CP 0 0.000045PF
C301_162 clk__L1_N0_426 0 0.000121PF
C302_162 clk__L1_N0_416 0 0.000625PF
C303_162 clk_r_REG31_S2:CP 0 0.000045PF
C304_162 clk__L1_N0_456 0 0.000121PF
C305_162 clk__L1_N0_451 0 0.000200PF
C306_162 clk__L1_N0_445 0 0.000219PF
C307_162 clk__L1_N0_436 0 0.000219PF
C308_162 clk__L1_N0_425 0 0.000518PF
C309_162 oDFF_12_q_reg:CP 0 0.000045PF
C310_162 clk__L1_N0_470 0 0.000121PF
C311_162 clk__L1_N0_466 0 0.000070PF
C312_162 clk__L1_N0_463 0 0.000426PF
C313_162 clk__L1_N0_459 0 0.000299PF
C314_162 clk__L1_N0_455 0 0.000184PF
C315_162 iDFF_14_q_reg:CP 0 0.000045PF
C316_162 clk__L1_N0_472 0 0.000121PF
C317_162 clk__L1_N0_469 0 0.000070PF
C318_162 oDFF_10_q_reg:CP 0 0.000045PF
C319_162 clk__L1_N0_477 0 0.000146PF
C320_162 clk__L1_N0_476 0 0.000306PF
C321_162 clk__L1_I0:Z 0 0.000435PF
C322_162 clk__L1_N0_471 0 0.000121PF
C323_162 clk__L1_N0_468 0 0.000121PF
C324_162 clk__L1_N0_465 0 0.000146PF
C325_162 clk_r_REG33_S2:CP 0 0.000045PF
C326_162 clk__L1_N0_496 0 0.000121PF
C327_162 clk__L1_N0_492 0 0.000130PF
C328_162 clk__L1_N0_489 0 0.000130PF
C329_162 clk__L1_N0_485 0 0.000371PF
C330_162 clk__L1_N0_482 0 0.000245PF
C331_162 clk__L1_N0_480 0 0.000204PF
C332_162 clk__L1_N0_478 0 0.000046PF
C333_162 clk_r_REG19_S2:CP 0 0.000045PF
C334_162 clk__L1_N0_495 0 0.000121PF
C335_162 clk__L1_N0_491 0 0.000410PF
C336_162 clk__L1_N0_488 0 0.000145PF
C337_162 clk_r_REG20_S2:CP 0 0.000045PF
C338_162 clk__L1_N0_499 0 0.000121PF
C339_162 clk__L1_N0_494 0 0.000394PF
C340_162 oDFF_14_q_reg:CP 0 0.000045PF
C341_162 clk__L1_N0_484 0 0.000121PF
C342_162 clk__L1_N0_481 0 0.000177PF
C343_162 iDFF_11_q_reg:CP 0 0.000045PF
C344_162 clk__L1_N0_498 0 0.000121PF
C345_162 clk__L1_N0_493 0 0.000235PF
C346_162 clk__L1_N0_490 0 0.000097PF
C347_162 clk__L1_N0_486 0 0.000153PF
C348_162 clk__L1_N0_483 0 0.000153PF
C349_162 clk_r_REG30_S2:CP 0 0.000045PF
C350_162 clk__L1_N0_504 0 0.000121PF
C351_162 clk__L1_N0_497 0 0.000413PF
C352_162 iDFF_15_q_reg:CP 0 0.000045PF
C353_162 clk__L1_N0_514 0 0.000121PF
C354_162 clk__L1_N0_512 0 0.000062PF
C355_162 clk__L1_N0_511 0 0.000062PF
C356_162 clk__L1_N0_508 0 0.000153PF
C357_162 clk__L1_N0_503 0 0.000153PF
C358_162 clk_r_REG34_S2:CP 0 0.000045PF
C359_162 clk__L1_N0_521 0 0.000121PF
C360_162 clk__L1_N0_518 0 0.000121PF
C361_162 clk__L1_N0_515 0 0.000324PF
C362_162 clk__L1_N0_513 0 0.000194PF
C363_162 clk_r_REG9_S2:CP 0 0.000045PF
C364_162 clk__L1_N0_530 0 0.000121PF
C365_162 clk__L1_N0_524 0 0.000398PF
C366_162 clk__L1_N0_520 0 0.000302PF
C367_162 clk__L1_N0_517 0 0.000324PF
C368_162 iDFF_3_q_reg:CP 0 0.000045PF
C369_162 clk__L1_N0_556 0 0.000121PF
C370_162 clk__L1_N0_549 0 0.000121PF
C371_162 clk__L1_N0_542 0 0.000194PF
C372_162 clk__L1_N0_535 0 0.000194PF
C373_162 clk__L1_N0_529 0 0.000254PF
C374_162 oDFF_15_q_reg:CP 0 0.000045PF
C375_162 clk__L1_N0_565 0 0.000121PF
C376_162 clk__L1_N0_560 0 0.000045PF
C377_162 clk__L1_N0_555 0 0.000045PF
C378_162 clk__L1_N0_548 0 0.000321PF
C379_162 clk__L1_N0_541 0 0.000321PF
C380_162 clk__L1_N0_534 0 0.000202PF
C381_162 oDFF_2_q_reg:CP 0 0.000045PF
C382_162 clk__L1_N0_554 0 0.000121PF
C383_162 clk__L1_N0_547 0 0.000089PF
C384_162 clk__L1_N0_540 0 0.000123PF
C385_162 iDFF_2_q_reg:CP 0 0.000045PF
C386_162 clk__L1_N0_528 0 0.000121PF
C387_162 clk__L1_N0_523 0 0.000121PF
C388_162 clk__L1_N0_519 0 0.000504PF
C389_162 clk_r_REG10_S2:CP 0 0.000045PF
C390_162 clk__L1_N0_564 0 0.000121PF
C391_162 clk__L1_N0_558 0 0.000053PF
C392_162 clk__L1_N0_553 0 0.000053PF
C393_162 clk__L1_N0_546 0 0.000208PF
C394_162 clk__L1_N0_539 0 0.000208PF
C395_162 clk__L1_N0_532 0 0.000351PF
C396_162 clk__L1_N0_527 0 0.000307PF
C397_162 clk__L1_N0_522 0 0.000457PF
C398_162 clk_r_REG5_S2:CP 0 0.000045PF
C399_162 clk__L1_N0_545 0 0.000121PF
C400_162 clk__L1_N0_538 0 0.000274PF
C401_162 oDFF_7_q_reg:CP 0 0.000045PF
C402_162 clk__L1_N0_563 0 0.000121PF
C403_162 clk__L1_N0_557 0 0.000060PF
C404_162 clk__L1_N0_551 0 0.000095PF
C405_162 clk__L1_N0_544 0 0.000264PF
C406_162 iDFF_7_q_reg:CP 0 0.000045PF
C407_162 clk__L1_N0_575 0 0.000121PF
C408_162 clk__L1_N0_573 0 0.000129PF
C409_162 clk__L1_N0_571 0 0.000129PF
C410_162 clk__L1_N0_566 0 0.000330PF
C411_162 clk__L1_N0_562 0 0.000213PF
C412_162 oDFF_3_q_reg:CP 0 0.000045PF
C413_162 clk__L1_N0_574 0 0.000121PF
C414_162 clk__L1_N0_572 0 0.000121PF
C415_162 clk__L1_N0_570 0 0.000136PF
C416_162 iDFF_6_q_reg:CP 0 0.000045PF
C417_162 clk__L1_N0_543 0 0.000121PF
C418_162 clk__L1_N0_537 0 0.000071PF
C419_162 clk__L1_N0_531 0 0.000071PF
C420_162 clk__L1_N0_526 0 0.000148PF
C421_162 oDFF_11_q_reg:CP 0 0.000045PF
C422_162 clk__L1_N0_507 0 0.000121PF
C423_162 clk__L1_N0_502 0 0.000276PF
C424_162 iDFF_10_q_reg:CP 0 0.000045PF
C425_162 clk__L1_N0_458 0 0.000121PF
C426_162 clk__L1_N0_454 0 0.000121PF
C427_162 clk__L1_N0_450 0 0.000878PF
C428_162 clk__L1_N0_444 0 0.000287PF
C429_162 clk__L1_N0_435 0 0.000333PF
C430_162 iDFF_36_q_reg:CP 0 0.000045PF
C431_162 clk__L1_N0_464 0 0.000121PF
C432_162 clk__L1_N0_461 0 0.000257PF
C433_162 clk__L1_N0_457 0 0.000257PF
C434_162 clk__L1_N0_453 0 0.000610PF
C435_162 clk_r_REG29_S2:CP 0 0.000045PF
C436_162 clk__L1_N0_449 0 0.000121PF
C437_162 clk__L1_N0_443 0 0.000132PF
C438_162 clk_r_REG32_S2:CP 0 0.000045PF
C439_162 clk__L1_N0_361 0 0.000033PF
C440_162 clk__L1_N0_351 0 0.000050PF
C441_162 clk__L1_N0_343 0 0.000297PF
C442_162 oDFF_16_q_reg:CP 0 0.000045PF
C443_162 clk__L1_N0_371 0 0.000035PF
C444_162 clk__L1_N0_360 0 0.000051PF
C445_162 clk__L1_N0_350 0 0.000387PF
C446_162 clk_r_REG35_S2:CP 0 0.000045PF
C447_162 clk__L1_N0_394 0 0.000121PF
C448_162 clk__L1_N0_382 0 0.000165PF
C449_162 clk__L1_N0_370 0 0.000091PF
C450_162 clk__L1_N0_359 0 0.000229PF
C451_162 iDFF_16_q_reg:CP 0 0.000045PF
C452_162 clk__L1_N0_404 0 0.000121PF
C453_162 clk__L1_N0_393 0 0.000127PF
C454_162 iDFF_4_q_reg:CP 0 0.000045PF
C455_162 clk__L1_N0_304 0 0.000121PF
C456_162 clk__L1_N0_299 0 0.000121PF
C457_162 clk__L1_N0_294 0 0.000189PF
C458_162 clk__L1_N0_289 0 0.000189PF
C459_162 clk__L1_N0_282 0 0.000164PF
C460_162 clk_r_REG22_S2:CP 0 0.000045PF
C461_162 clk__L1_N0_212 0 0.000121PF
C462_162 clk__L1_N0_205 0 0.000459PF
C463_162 clk_r_REG3_S2:CP 0 0.000045PF
C464_162 clk__L1_N0_217 0 0.000121PF
C465_162 clk__L1_N0_211 0 0.000352PF
C466_162 clk_r_REG17_S2:CP 0 0.000045PF
C467_162 clk__L1_N0_246 0 0.000121PF
C468_162 clk__L1_N0_240 0 0.000399PF
C469_162 clk__L1_N0_232 0 0.000092PF
C470_162 clk__L1_N0_224 0 0.000189PF
C471_162 clk__L1_N0_216 0 0.000189PF
C472_162 clk_r_REG4_S2:CP 0 0.000045PF
C473_162 clk__L1_N0_273 0 0.000121PF
C474_162 clk__L1_N0_266 0 0.000261PF
C475_162 clk__L1_N0_260 0 0.000103PF
C476_162 clk__L1_N0_252 0 0.000103PF
C477_162 clk__L1_N0_245 0 0.000345PF
C478_162 iDFF_33_q_reg:CP 0 0.000045PF
C479_162 clk__L1_N0_308 0 0.000067PF
C480_162 clk__L1_N0_303 0 0.000067PF
C481_162 clk__L1_N0_298 0 0.000166PF
C482_162 clk__L1_N0_293 0 0.000166PF
C483_162 clk__L1_N0_288 0 0.000147PF
C484_162 clk__L1_N0_280 0 0.000331PF
C485_162 clk__L1_N0_272 0 0.000245PF
C486_162 iDFF_34_q_reg:CP 0 0.000045PF
C487_162 clk__L1_N0_319 0 0.000121PF
C488_162 clk__L1_N0_316 0 0.000766PF
C489_162 clk__L1_N0_313 0 0.000500PF
C490_162 iDFF_38_q_reg:CP 0 0.000045PF
C491_162 clk__L1_N0_342 0 0.000121PF
C492_162 clk__L1_N0_337 0 0.000121PF
C493_162 clk__L1_N0_330 0 0.000170PF
C494_162 clk__L1_N0_323 0 0.000170PF
C495_162 clk__L1_N0_318 0 0.000687PF
C496_162 iDFF_37_q_reg:CP 0 0.000045PF
C497_162 clk__L1_N0_329 0 0.000121PF
C498_162 clk__L1_N0_322 0 0.000421PF
C499_162 iDFF_41_q_reg:CP 0 0.000045PF
C500_162 clk__L1_N0_358 0 0.000121PF
C501_162 clk__L1_N0_348 0 0.000350PF
C502_162 clk__L1_N0_341 0 0.000093PF
C503_162 clk__L1_N0_335 0 0.000148PF
C504_162 clk__L1_N0_328 0 0.000148PF
C505_162 clk_r_REG13_S2:CP 0 0.000045PF
C506_162 clk__L1_N0_403 0 0.000121PF
C507_162 clk__L1_N0_392 0 0.000175PF
C508_162 clk__L1_N0_381 0 0.000175PF
C509_162 clk__L1_N0_368 0 0.000362PF
C510_162 clk__L1_N0_357 0 0.000362PF
C511_162 iDFF_18_q_reg:CP 0 0.000045PF
C512_162 clk__L1_N0_367 0 0.000121PF
C513_162 clk__L1_N0_356 0 0.000373PF
C514_162 clk_r_REG28_S2:CP 0 0.000045PF
C515_162 clk__L1_N0_413 0 0.000121PF
C516_162 clk__L1_N0_402 0 0.000121PF
C517_162 clk__L1_N0_391 0 0.000213PF
C518_162 clk__L1_N0_379 0 0.000213PF
C519_162 clk__L1_N0_366 0 0.000136PF
C520_162 clk_r_REG37_S2:CP 0 0.000045PF
C521_162 clk__L1_N0_390 0 0.000121PF
C522_162 clk__L1_N0_378 0 0.000640PF
C523_162 oDFF_18_q_reg:CP 0 0.000045PF
C524_162 clk__L1_N0_400 0 0.000121PF
C525_162 clk__L1_N0_389 0 0.000943PF
C526_162 clk_r_REG6_S2:CP 0 0.000045PF
C527_162 clk__L1_N0_434 0 0.000121PF
C528_162 clk__L1_N0_423 0 0.000188PF
C529_162 clk__L1_N0_411 0 0.000148PF
C530_162 clk__L1_N0_399 0 0.000450PF
C531_162 iDFF_35_q_reg:CP 0 0.000045PF
C532_162 clk__L1_N0_441 0 0.000121PF
C533_162 clk__L1_N0_433 0 0.000188PF
C534_162 clk_r_REG41_S2:CP 0 0.000045PF
C535_162 clk__L1_N0_432 0 0.000121PF
C536_162 clk__L1_N0_422 0 0.000545PF
C537_162 clk__L1_N0_410 0 0.000321PF
C538_162 iDFF_22_q_reg:CP 0 0.000045PF
C539_162 clk__L1_N0_439 0 0.000121PF
C540_162 clk__L1_N0_431 0 0.000388PF
C541_162 iDFF_40_q_reg:CP 0 0.000045PF
C542_162 clk__L1_N0_438 0 0.000121PF
C543_162 clk__L1_N0_430 0 0.000176PF
C544_162 oDFF_22_q_reg:CP 0 0.000045PF
C545_162 clk__L1_N0_409 0 0.000086PF
C546_162 clk__L1_N0_398 0 0.000343PF
C547_162 oDFF_6_q_reg:CP 0 0.000045PF
C548_162 clk__L1_N0_420 0 0.000086PF
C549_162 iDFF_39_q_reg:CP 0 0.000045PF
C550_162 clk__L1_N0_297 0 0.000121PF
C551_162 clk__L1_N0_292 0 0.000121PF
C552_162 clk__L1_N0_287 0 0.000203PF
C553_162 clk_r_REG18_S2:CP 0 0.000045PF
C554_162 clk__L1_N0_259 0 0.000121PF
C555_162 clk__L1_N0_251 0 0.000038PF
C556_162 clk_r_REG21_S2:CP 0 0.000045PF
C557_162 clk__L1_N0_204 0 0.000121PF
C558_162 clk__L1_N0_198 0 0.000032PF
C559_162 oDFF_31_q_reg:CP 0 0.000045PF
C560_162 clk__L1_N0_68 0 0.000121PF
C561_162 clk__L1_N0_59 0 0.000760PF
C562_162 oDFF_32_q_reg:CP 0 0.000045PF
C563_162 clk__L1_N0_96 0 0.000121PF
C564_162 clk__L1_N0_90 0 0.000129PF
C565_162 clk__L1_N0_84 0 0.000129PF
C566_162 clk__L1_N0_76 0 0.000195PF
C567_162 clk__L1_N0_67 0 0.000195PF
C568_162 oDFF_25_q_reg:CP 0 0.000045PF
C569_162 clk__L1_N0_75 0 0.000121PF
C570_162 clk__L1_N0_66 0 0.000382PF
C571_162 clk_r_REG47_S2:CP 0 0.000045PF
C572_162 clk__L1_N0_19 0 0.000121PF
C573_162 clk__L1_N0_13 0 0.000117PF
C574_162 oDFF_23_q_reg:CP 0 0.000045PF
C575_162 clk__L1_N0_6 0 0.000121PF
C576_162 clk__L1_N0_3 0 0.000121PF
C577_162 clk__L1_N0_1 0 0.000090PF
R1_162 clk__L1_N0_2 clk__L1_N0_1 0.912000
R2_162 clk__L1_N0_1 clk__L1_N0_3 4.000000
R3_162 clk__L1_N0_4 clk__L1_N0_2 3.040000
R4_162 clk__L1_N0_2 clk__L1_N0_5 4.000000
R5_162 clk__L1_N0_3 clk__L1_N0_6 4.000000
R6_162 clk__L1_N0_4 clk__L1_N0_7 4.000000
R7_162 clk__L1_N0_5 clk__L1_N0_8 3.344000
R8_162 clk__L1_N0_6 oDFF_23_q_reg:CP 4.000000
R9_162 clk__L1_N0_10 clk__L1_N0_7 5.016000
R10_162 clk__L1_N0_7 clk__L1_N0_11 1.672000
R11_162 clk__L1_N0_8 clk__L1_N0_12 4.000000
R12_162 clk__L1_N0_13 clk__L1_N0_10 0.912000
R13_162 clk__L1_N0_10 clk__L1_N0_14 4.000000
R14_162 clk__L1_N0_10 clk__L1_N0_15 4.000000
R15_162 clk__L1_N0_11 clk__L1_N0_16 2.736000
R16_162 clk__L1_N0_11 clk__L1_N0_17 4.000000
R17_162 clk__L1_N0_18 clk__L1_N0_12 1.368000
R18_162 clk__L1_N0_13 clk__L1_N0_19 4.000000
R19_162 clk__L1_N0_14 clk__L1_N0_20 1.672000
R20_162 clk__L1_N0_15 iDFF_28_q_reg:CP 4.000000
R21_162 clk__L1_N0_16 clk__L1_N0_22 3.496000
R22_162 clk__L1_N0_16 clk__L1_N0_23 4.000000
R23_162 clk__L1_N0_17 oDFF_19_q_reg:CP 4.000000
R24_162 clk__L1_N0_18 clk__L1_N0_25 4.000000
R25_162 clk__L1_N0_19 clk_r_REG47_S2:CP 4.000000
R26_162 clk__L1_N0_20 clk__L1_N0_27 4.000000
R27_162 clk__L1_N0_22 clk__L1_N0_28 6.992000
R28_162 clk__L1_N0_22 clk__L1_N0_29 4.000000
R29_162 clk__L1_N0_30 clk__L1_N0_23 2.280000
R30_162 clk__L1_N0_25 clk__L1_N0_31 0.608000
R31_162 clk__L1_N0_25 clk__L1_N0_32 4.000000
R32_162 clk__L1_N0_33 clk__L1_N0_27 2.584000
R33_162 clk__L1_N0_27 clk__L1_N0_34 4.000000
R34_162 clk__L1_N0_28 clk__L1_N0_35 4.000000
R35_162 clk__L1_N0_28 clk__L1_N0_36 4.000000
R36_162 clk__L1_N0_29 clk_r_REG39_S2:CP 4.000000
R37_162 clk__L1_N0_30 clk__L1_N0_38 4.000000
R38_162 clk__L1_N0_31 clk__L1_N0_39 2.280000
R39_162 clk__L1_N0_31 clk__L1_N0_40 4.000000
R40_162 clk__L1_N0_32 clk_r_REG42_S2:CP 4.000000
R41_162 clk__L1_N0_42 clk__L1_N0_33 0.912000
R42_162 clk__L1_N0_33 clk__L1_N0_43 4.000000
R43_162 clk__L1_N0_34 iDFF_32_q_reg:CP 4.000000
R44_162 clk__L1_N0_45 clk__L1_N0_35 2.280000
R45_162 clk__L1_N0_36 clk_r_REG43_S2:CP 4.000000
R46_162 clk__L1_N0_38 clk__L1_N0_47 4.000000
R47_162 clk__L1_N0_39 clk__L1_N0_48 4.408000
R48_162 clk__L1_N0_39 clk__L1_N0_49 4.000000
R49_162 clk__L1_N0_40 iDFF_23_q_reg:CP 4.000000
R50_162 clk__L1_N0_51 clk__L1_N0_42 2.432000
R51_162 clk__L1_N0_42 clk__L1_N0_52 4.000000
R52_162 clk__L1_N0_43 iDFF_31_q_reg:CP 4.000000
R53_162 clk__L1_N0_45 clk__L1_N0_54 4.000000
R54_162 clk__L1_N0_47 clk_r_REG38_S2:CP 4.000000
R55_162 clk__L1_N0_48 clk__L1_N0_56 5.320000
R56_162 clk__L1_N0_48 clk__L1_N0_57 4.000000
R57_162 clk__L1_N0_49 iDFF_20_q_reg:CP 4.000000
R58_162 clk__L1_N0_59 clk__L1_N0_51 4.712000
R59_162 clk__L1_N0_51 clk__L1_N0_60 4.000000
R60_162 clk__L1_N0_51 clk__L1_N0_61 4.000000
R61_162 clk__L1_N0_52 oDFF_28_q_reg:CP 4.000000
R62_162 clk__L1_N0_54 clk__L1_N0_63 0.456000
R63_162 clk__L1_N0_56 clk__L1_N0_64 4.000000
R64_162 clk__L1_N0_57 clk__L1_N0_65 2.280000
R65_162 clk__L1_N0_66 clk__L1_N0_59 4.712000
R66_162 clk__L1_N0_59 clk__L1_N0_67 4.000000
R67_162 clk__L1_N0_59 clk__L1_N0_68 4.000000
R68_162 clk__L1_N0_69 clk__L1_N0_60 1.672000
R69_162 clk__L1_N0_61 clk_r_REG51_S2:CP 4.000000
R70_162 clk__L1_N0_63 clk__L1_N0_71 4.000000
R71_162 clk__L1_N0_63 clk__L1_N0_72 4.000000
R72_162 clk__L1_N0_64 iDFF_24_q_reg:CP 4.000000
R73_162 clk__L1_N0_65 clk__L1_N0_74 4.000000
R74_162 clk__L1_N0_66 clk__L1_N0_75 4.000000
R75_162 clk__L1_N0_67 clk__L1_N0_76 2.280000
R76_162 clk__L1_N0_68 oDFF_31_q_reg:CP 4.000000
R77_162 clk__L1_N0_78 clk__L1_N0_69 2.280000
R78_162 clk__L1_N0_69 clk__L1_N0_79 4.000000
R79_162 clk__L1_N0_80 clk__L1_N0_71 1.672000
R80_162 clk__L1_N0_72 oDFF_24_q_reg:CP 4.000000
R81_162 clk__L1_N0_74 clk__L1_N0_82 4.000000
R82_162 clk__L1_N0_75 oDFF_25_q_reg:CP 4.000000
R83_162 clk__L1_N0_76 clk__L1_N0_84 4.000000
R84_162 clk__L1_N0_85 clk__L1_N0_78 1.520000
R85_162 clk__L1_N0_78 clk__L1_N0_86 4.000000
R86_162 clk__L1_N0_79 clk__L1_N0_87 0.304000
R87_162 clk__L1_N0_80 clk__L1_N0_88 4.000000
R88_162 clk__L1_N0_82 oDFF_20_q_reg:CP 4.000000
R89_162 clk__L1_N0_84 clk__L1_N0_90 1.368000
R90_162 clk__L1_N0_85 clk__L1_N0_91 4.000000
R91_162 clk__L1_N0_86 clk__L1_N0_92 2.432000
R92_162 clk__L1_N0_86 clk__L1_N0_93 4.000000
R93_162 clk__L1_N0_87 clk__L1_N0_94 4.000000
R94_162 clk__L1_N0_88 clk__L1_N0_95 1.672000
R95_162 clk__L1_N0_90 clk__L1_N0_96 4.000000
R96_162 clk__L1_N0_97 clk__L1_N0_91 2.888000
R97_162 clk__L1_N0_92 clk__L1_N0_98 4.000000
R98_162 clk__L1_N0_92 clk__L1_N0_99 4.000000
R99_162 clk__L1_N0_93 oDFF_27_q_reg:CP 4.000000
R100_162 clk__L1_N0_94 clk_r_REG50_S2:CP 4.000000
R101_162 clk__L1_N0_95 clk__L1_N0_102 4.000000
R102_162 clk__L1_N0_96 oDFF_32_q_reg:CP 4.000000
R103_162 clk__L1_N0_97 clk__L1_N0_104 4.000000
R104_162 clk__L1_N0_97 clk__L1_N0_105 4.000000
R105_162 clk__L1_N0_106 clk__L1_N0_98 1.672000
R106_162 clk__L1_N0_99 clk_r_REG44_S2:CP 4.000000
R107_162 clk__L1_N0_102 iDFF_21_q_reg:CP 4.000000
R108_162 clk__L1_N0_109 clk__L1_N0_104 2.432000
R109_162 clk__L1_N0_105 clk_r_REG24_S2:CP 4.000000
R110_162 clk__L1_N0_106 clk__L1_N0_111 4.000000
R111_162 clk__L1_N0_109 clk__L1_N0_112 0.152000
R112_162 clk__L1_N0_109 clk__L1_N0_113 4.000000
R113_162 clk__L1_N0_114 clk__L1_N0_111 0.152000
R114_162 clk__L1_N0_111 clk__L1_N0_115 0.912000
R115_162 clk__L1_N0_116 clk__L1_N0_112 1.368000
R116_162 clk__L1_N0_117 clk__L1_N0_113 2.128000
R117_162 clk__L1_N0_113 clk__L1_N0_118 0.304000
R118_162 clk__L1_N0_114 clk__L1_N0_119 4.000000
R119_162 clk__L1_N0_115 clk__L1_N0_120 4.000000
R120_162 clk__L1_N0_115 clk__L1_N0_121 4.000000
R121_162 clk__L1_N0_122 clk__L1_N0_116 2.584000
R122_162 clk__L1_N0_116 clk__L1_N0_123 4.000000
R123_162 clk__L1_N0_124 clk__L1_N0_117 4.104000
R124_162 clk__L1_N0_117 clk__L1_N0_125 4.000000
R125_162 clk__L1_N0_118 clk__L1_N0_126 4.000000
R126_162 clk__L1_N0_119 clk_r_REG46_S2:CP 4.000000
R127_162 clk__L1_N0_128 clk__L1_N0_120 2.128000
R128_162 clk__L1_N0_121 iDFF_27_q_reg:CP 4.000000
R129_162 clk__L1_N0_130 clk__L1_N0_122 1.672000
R130_162 clk__L1_N0_122 clk__L1_N0_131 4.000000
R131_162 clk__L1_N0_123 clk__L1_N0_132 4.000000
R132_162 clk__L1_N0_133 clk__L1_N0_124 0.760000
R133_162 clk__L1_N0_124 clk__L1_N0_134 4.000000
R134_162 clk__L1_N0_124 clk__L1_N0_135 4.000000
R135_162 clk__L1_N0_125 clk__L1_N0_136 0.152000
R136_162 clk__L1_N0_126 clk_r_REG15_S2:CP 4.000000
R137_162 clk__L1_N0_128 clk__L1_N0_138 4.000000
R138_162 clk__L1_N0_130 clk__L1_N0_139 4.000000
R139_162 clk__L1_N0_131 clk__L1_N0_140 0.152000
R140_162 clk__L1_N0_141 clk__L1_N0_132 0.304000
R141_162 clk__L1_N0_142 clk__L1_N0_133 1.368000
R142_162 clk__L1_N0_133 clk__L1_N0_143 4.000000
R143_162 clk__L1_N0_134 clk__L1_N0_144 2.280000
R144_162 clk__L1_N0_145 clk__L1_N0_134 1.672000
R145_162 clk__L1_N0_135 iDFF_26_q_reg:CP 4.000000
R146_162 clk__L1_N0_136 clk_r_REG12_S2:CP 4.000000
R147_162 clk__L1_N0_138 clk__L1_N0_148 0.456000
R148_162 clk__L1_N0_149 clk__L1_N0_139 1.976000
R149_162 clk__L1_N0_140 clk__L1_N0_150 4.000000
R150_162 clk__L1_N0_141 clk_r_REG45_S2:CP 4.000000
R151_162 clk__L1_N0_152 clk__L1_N0_142 0.304000
R152_162 clk__L1_N0_142 clk__L1_N0_153 4.000000
R153_162 clk__L1_N0_143 oDFF_26_q_reg:CP 4.000000
R154_162 clk__L1_N0_144 clk__L1_N0_155 4.000000
R155_162 clk__L1_N0_145 clk__L1_N0_156 4.000000
R156_162 clk__L1_N0_148 clk__L1_N0_157 4.104000
R157_162 clk__L1_N0_148 clk__L1_N0_158 4.000000
R158_162 clk__L1_N0_159 clk__L1_N0_149 5.016000
R159_162 clk__L1_N0_149 clk__L1_N0_160 4.000000
R160_162 clk__L1_N0_150 clk_r_REG27_S2:CP 4.000000
R161_162 clk__L1_N0_152 clk__L1_N0_162 4.000000
R162_162 clk__L1_N0_153 clk__L1_N0_163 3.952000
R163_162 clk__L1_N0_155 clk__L1_N0_164 0.760000
R164_162 clk__L1_N0_156 clk__L1_N0_165 1.672000
R165_162 clk__L1_N0_166 clk__L1_N0_157 0.152000
R166_162 clk__L1_N0_158 clk_r_REG16_S2:CP 4.000000
R167_162 clk__L1_N0_159 clk__L1_N0_168 4.000000
R168_162 clk__L1_N0_159 clk__L1_N0_169 4.000000
R169_162 clk__L1_N0_160 clk_r_REG14_S2:CP 4.000000
R170_162 clk__L1_N0_171 clk__L1_N0_162 1.672000
R171_162 clk__L1_N0_163 clk__L1_N0_172 4.000000
R172_162 clk__L1_N0_164 clk__L1_N0_173 4.000000
R173_162 clk__L1_N0_165 clk__L1_N0_174 4.000000
R174_162 clk__L1_N0_166 clk__L1_N0_175 0.456000
R175_162 clk__L1_N0_176 clk__L1_N0_168 2.280000
R176_162 clk__L1_N0_169 oDFF_30_q_reg:CP 4.000000
R177_162 clk__L1_N0_171 clk__L1_N0_178 4.000000
R178_162 clk__L1_N0_172 clk__L1_N0_179 4.000000
R179_162 clk__L1_N0_173 clk_r_REG48_S2:CP 4.000000
R180_162 clk__L1_N0_174 clk_r_REG49_S2:CP 4.000000
R181_162 clk__L1_N0_175 clk__L1_N0_182 1.368000
R182_162 clk__L1_N0_175 clk__L1_N0_183 4.000000
R183_162 clk__L1_N0_184 clk__L1_N0_176 3.952000
R184_162 clk__L1_N0_176 clk__L1_N0_185 4.000000
R185_162 clk__L1_N0_178 clk__L1_N0_186 4.000000
R186_162 clk__L1_N0_179 oDFF_29_q_reg:CP 4.000000
R187_162 clk__L1_N0_182 clk__L1_N0_188 5.928000
R188_162 clk__L1_N0_182 clk__L1_N0_189 4.000000
R189_162 clk__L1_N0_190 clk__L1_N0_183 1.672000
R190_162 clk__L1_N0_184 clk__L1_N0_191 4.000000
R191_162 clk__L1_N0_185 clk__L1_N0_192 1.216000
R192_162 clk__L1_N0_186 iDFF_30_q_reg:CP 4.000000
R193_162 clk__L1_N0_188 clk__L1_N0_194 4.000000
R194_162 clk__L1_N0_188 clk__L1_N0_195 4.000000
R195_162 clk__L1_N0_189 iDFF_25_q_reg:CP 4.000000
R196_162 clk__L1_N0_190 clk__L1_N0_197 4.000000
R197_162 clk__L1_N0_198 clk__L1_N0_191 0.152000
R198_162 clk__L1_N0_191 clk__L1_N0_199 1.368000
R199_162 clk__L1_N0_192 clk__L1_N0_200 4.000000
R200_162 clk__L1_N0_194 clk__L1_N0_201 2.280000
R201_162 clk__L1_N0_195 iDFF_17_q_reg:CP 4.000000
R202_162 clk__L1_N0_197 clk__L1_N0_203 4.000000
R203_162 clk__L1_N0_198 clk__L1_N0_204 4.000000
R204_162 clk__L1_N0_199 clk__L1_N0_205 0.912000
R205_162 clk__L1_N0_199 clk__L1_N0_206 4.000000
R206_162 clk__L1_N0_200 clk_r_REG11_S2:CP 4.000000
R207_162 clk__L1_N0_201 clk__L1_N0_208 4.000000
R208_162 clk__L1_N0_203 iDFF_29_q_reg:CP 4.000000
R209_162 clk__L1_N0_204 clk_r_REG21_S2:CP 4.000000
R210_162 clk__L1_N0_205 clk__L1_N0_211 3.800000
R211_162 clk__L1_N0_205 clk__L1_N0_212 4.000000
R212_162 clk__L1_N0_213 clk__L1_N0_206 1.672000
R213_162 clk__L1_N0_208 clk__L1_N0_214 2.888000
R214_162 clk__L1_N0_208 clk__L1_N0_215 4.000000
R215_162 clk__L1_N0_211 clk__L1_N0_216 4.000000
R216_162 clk__L1_N0_211 clk__L1_N0_217 4.000000
R217_162 clk__L1_N0_212 clk_r_REG22_S2:CP 4.000000
R218_162 clk__L1_N0_213 clk__L1_N0_219 4.000000
R219_162 clk__L1_N0_214 clk__L1_N0_220 2.432000
R220_162 clk__L1_N0_214 clk__L1_N0_221 4.000000
R221_162 clk__L1_N0_214 clk__L1_N0_222 4.000000
R222_162 clk__L1_N0_215 iDFF_19_q_reg:CP 4.000000
R223_162 clk__L1_N0_216 clk__L1_N0_224 2.280000
R224_162 clk__L1_N0_217 clk_r_REG3_S2:CP 4.000000
R225_162 clk__L1_N0_226 clk__L1_N0_219 1.368000
R226_162 clk__L1_N0_219 clk__L1_N0_227 4.000000
R227_162 clk__L1_N0_220 clk__L1_N0_228 2.584000
R228_162 clk__L1_N0_220 clk__L1_N0_229 4.000000
R229_162 clk__L1_N0_230 clk__L1_N0_221 2.280000
R230_162 clk__L1_N0_222 clk__L1_N0_231 0.152000
R231_162 clk__L1_N0_224 clk__L1_N0_232 4.000000
R232_162 clk__L1_N0_226 clk__L1_N0_233 4.000000
R233_162 clk__L1_N0_227 clk_r_REG8_S2:CP 4.000000
R234_162 clk__L1_N0_228 clk__L1_N0_235 1.824000
R235_162 clk__L1_N0_228 clk__L1_N0_236 4.000000
R236_162 clk__L1_N0_229 clk_r_REG40_S2:CP 4.000000
R237_162 clk__L1_N0_230 clk__L1_N0_238 4.000000
R238_162 clk__L1_N0_231 clk_r_REG25_S2:CP 4.000000
R239_162 clk__L1_N0_232 clk__L1_N0_240 0.608000
R240_162 clk__L1_N0_241 clk__L1_N0_233 2.128000
R241_162 clk__L1_N0_235 clk__L1_N0_242 4.000000
R242_162 clk__L1_N0_236 oDFF_17_q_reg:CP 4.000000
R243_162 clk__L1_N0_238 clk__L1_N0_244 0.304000
R244_162 clk__L1_N0_240 clk__L1_N0_245 3.496000
R245_162 clk__L1_N0_240 clk__L1_N0_246 4.000000
R246_162 clk__L1_N0_247 clk__L1_N0_241 1.824000
R247_162 clk__L1_N0_241 clk__L1_N0_248 4.000000
R248_162 clk__L1_N0_249 clk__L1_N0_242 3.952000
R249_162 clk__L1_N0_244 clk__L1_N0_250 4.000000
R250_162 clk__L1_N0_245 clk__L1_N0_251 0.152000
R251_162 clk__L1_N0_245 clk__L1_N0_252 4.000000
R252_162 clk__L1_N0_246 clk_r_REG17_S2:CP 4.000000
R253_162 clk__L1_N0_254 clk__L1_N0_247 2.128000
R254_162 clk__L1_N0_247 clk__L1_N0_255 4.000000
R255_162 clk__L1_N0_248 clk__L1_N0_256 4.000000
R256_162 clk__L1_N0_249 clk__L1_N0_257 4.000000
R257_162 clk__L1_N0_250 clk_r_REG36_S2:CP 4.000000
R258_162 clk__L1_N0_251 clk__L1_N0_259 4.000000
R259_162 clk__L1_N0_252 clk__L1_N0_260 1.672000
R260_162 clk__L1_N0_254 clk__L1_N0_261 4.000000
R261_162 clk__L1_N0_255 clk__L1_N0_262 2.280000
R262_162 clk__L1_N0_256 oDFF_4_q_reg:CP 4.000000
R263_162 clk__L1_N0_257 clk__L1_N0_264 0.912000
R264_162 clk__L1_N0_259 clk_r_REG18_S2:CP 4.000000
R265_162 clk__L1_N0_260 clk__L1_N0_266 4.000000
R266_162 clk__L1_N0_267 clk__L1_N0_261 0.152000
R267_162 clk__L1_N0_261 clk__L1_N0_268 0.608000
R268_162 clk__L1_N0_262 clk__L1_N0_269 1.064000
R269_162 clk__L1_N0_262 clk__L1_N0_270 4.000000
R270_162 clk__L1_N0_264 clk__L1_N0_271 4.000000
R271_162 clk__L1_N0_266 clk__L1_N0_272 2.888000
R272_162 clk__L1_N0_266 clk__L1_N0_273 4.000000
R273_162 clk__L1_N0_274 clk__L1_N0_267 0.456000
R274_162 clk__L1_N0_267 clk__L1_N0_275 4.000000
R275_162 clk__L1_N0_268 clk__L1_N0_276 4.000000
R276_162 clk__L1_N0_269 clk__L1_N0_277 4.000000
R277_162 clk__L1_N0_270 clk_r_REG1_S2:CP 4.000000
R278_162 clk__L1_N0_271 oDFF_21_q_reg:CP 4.000000
R279_162 clk__L1_N0_272 clk__L1_N0_280 4.000000
R280_162 clk__L1_N0_273 clk_r_REG4_S2:CP 4.000000
R281_162 clk__L1_N0_282 clk__L1_N0_274 1.216000
R282_162 clk__L1_N0_274 clk__L1_N0_283 4.000000
R283_162 clk__L1_N0_275 oDFF_1_q_reg:CP 4.000000
R284_162 clk__L1_N0_285 clk__L1_N0_276 0.152000
R285_162 clk__L1_N0_277 iDFF_1_q_reg:CP 4.000000
R286_162 clk__L1_N0_280 clk__L1_N0_287 2.280000
R287_162 clk__L1_N0_288 clk__L1_N0_280 1.368000
R288_162 clk__L1_N0_282 clk__L1_N0_289 4.000000
R289_162 clk__L1_N0_290 clk__L1_N0_283 1.824000
R290_162 clk__L1_N0_285 iDFF_8_q_reg:CP 4.000000
R291_162 clk__L1_N0_287 clk__L1_N0_292 4.000000
R292_162 clk__L1_N0_288 clk__L1_N0_293 4.000000
R293_162 clk__L1_N0_289 clk__L1_N0_294 2.128000
R294_162 clk__L1_N0_295 clk__L1_N0_290 2.128000
R295_162 clk__L1_N0_290 clk__L1_N0_296 4.000000
R296_162 clk__L1_N0_292 clk__L1_N0_297 4.000000
R297_162 clk__L1_N0_293 clk__L1_N0_298 1.672000
R298_162 clk__L1_N0_294 clk__L1_N0_299 4.000000
R299_162 clk__L1_N0_295 clk__L1_N0_300 4.000000
R300_162 clk__L1_N0_296 clk__L1_N0_301 0.760000
R301_162 clk__L1_N0_297 iDFF_39_q_reg:CP 4.000000
R302_162 clk__L1_N0_298 clk__L1_N0_303 4.000000
R303_162 clk__L1_N0_299 clk__L1_N0_304 4.000000
R304_162 clk__L1_N0_300 clk__L1_N0_305 2.128000
R305_162 clk__L1_N0_300 clk__L1_N0_306 4.000000
R306_162 clk__L1_N0_301 clk__L1_N0_307 4.000000
R307_162 clk__L1_N0_308 clk__L1_N0_303 0.304000
R308_162 clk__L1_N0_304 iDFF_4_q_reg:CP 4.000000
R309_162 clk__L1_N0_305 clk__L1_N0_310 4.000000
R310_162 clk__L1_N0_306 oDFF_8_q_reg:CP 4.000000
R311_162 clk__L1_N0_307 clk_r_REG7_S2:CP 4.000000
R312_162 clk__L1_N0_308 clk__L1_N0_313 4.000000
R313_162 clk__L1_N0_308 iDFF_33_q_reg:CP 4.000000
R314_162 clk__L1_N0_315 clk__L1_N0_310 1.672000
R315_162 clk__L1_N0_313 clk__L1_N0_316 3.800000
R316_162 clk__L1_N0_315 clk__L1_N0_317 4.000000
R317_162 clk__L1_N0_316 clk__L1_N0_318 1.976000
R318_162 clk__L1_N0_316 clk__L1_N0_319 4.000000
R319_162 clk__L1_N0_317 clk__L1_N0_320 2.280000
R320_162 clk__L1_N0_317 clk__L1_N0_321 4.000000
R321_162 clk__L1_N0_318 clk__L1_N0_322 4.104000
R322_162 clk__L1_N0_318 clk__L1_N0_323 4.000000
R323_162 clk__L1_N0_319 iDFF_34_q_reg:CP 4.000000
R324_162 clk__L1_N0_320 clk__L1_N0_325 1.368000
R325_162 clk__L1_N0_320 clk__L1_N0_326 4.000000
R326_162 clk__L1_N0_327 clk__L1_N0_321 0.152000
R327_162 clk__L1_N0_322 clk__L1_N0_328 4.000000
R328_162 clk__L1_N0_322 clk__L1_N0_329 4.000000
R329_162 clk__L1_N0_323 clk__L1_N0_330 1.672000
R330_162 clk__L1_N0_325 clk__L1_N0_331 2.584000
R331_162 clk__L1_N0_325 clk__L1_N0_332 4.000000
R332_162 clk__L1_N0_326 oDFF_5_q_reg:CP 4.000000
R333_162 clk__L1_N0_327 clk_r_REG2_S2:CP 4.000000
R334_162 clk__L1_N0_328 clk__L1_N0_335 1.672000
R335_162 clk__L1_N0_329 iDFF_37_q_reg:CP 4.000000
R336_162 clk__L1_N0_330 clk__L1_N0_337 4.000000
R337_162 clk__L1_N0_331 clk__L1_N0_338 2.432000
R338_162 clk__L1_N0_331 clk__L1_N0_339 4.000000
R339_162 clk__L1_N0_332 clk__L1_N0_340 1.520000
R340_162 clk__L1_N0_335 clk__L1_N0_341 4.000000
R341_162 clk__L1_N0_337 clk__L1_N0_342 4.000000
R342_162 clk__L1_N0_338 clk__L1_N0_343 1.064000
R343_162 clk__L1_N0_338 clk__L1_N0_344 4.000000
R344_162 clk__L1_N0_345 clk__L1_N0_339 0.152000
R345_162 clk__L1_N0_340 clk__L1_N0_346 2.432000
R346_162 clk__L1_N0_340 clk__L1_N0_347 4.000000
R347_162 clk__L1_N0_341 clk__L1_N0_348 0.608000
R348_162 clk__L1_N0_342 iDFF_38_q_reg:CP 4.000000
R349_162 clk__L1_N0_343 clk__L1_N0_350 2.280000
R350_162 clk__L1_N0_343 clk__L1_N0_351 4.000000
R351_162 clk__L1_N0_344 clk__L1_N0_352 1.520000
R352_162 clk__L1_N0_345 oDFF_13_q_reg:CP 4.000000
R353_162 clk__L1_N0_346 clk__L1_N0_354 4.000000
R354_162 clk__L1_N0_347 clk__L1_N0_355 4.000000
R355_162 clk__L1_N0_348 clk__L1_N0_356 2.280000
R356_162 clk__L1_N0_348 clk__L1_N0_357 4.000000
R357_162 clk__L1_N0_348 clk__L1_N0_358 4.000000
R358_162 clk__L1_N0_350 clk__L1_N0_359 1.824000
R359_162 clk__L1_N0_350 clk__L1_N0_360 4.000000
R360_162 clk__L1_N0_361 clk__L1_N0_351 0.152000
R361_162 clk__L1_N0_352 clk__L1_N0_362 2.280000
R362_162 clk__L1_N0_352 clk__L1_N0_363 4.000000
R363_162 clk__L1_N0_354 clk__L1_N0_364 0.304000
R364_162 clk__L1_N0_355 iDFF_5_q_reg:CP 4.000000
R365_162 clk__L1_N0_356 clk__L1_N0_366 0.912000
R366_162 clk__L1_N0_356 clk__L1_N0_367 4.000000
R367_162 clk__L1_N0_357 clk__L1_N0_368 4.104000
R368_162 clk__L1_N0_358 iDFF_41_q_reg:CP 4.000000
R369_162 clk__L1_N0_370 clk__L1_N0_359 0.152000
R370_162 clk__L1_N0_371 clk__L1_N0_360 0.152000
R371_162 clk__L1_N0_361 clk_r_REG32_S2:CP 4.000000
R372_162 clk__L1_N0_362 clk__L1_N0_373 1.672000
R373_162 clk__L1_N0_362 clk__L1_N0_374 4.000000
R374_162 clk__L1_N0_363 clk__L1_N0_375 4.000000
R375_162 clk__L1_N0_364 clk__L1_N0_376 1.368000
R376_162 clk__L1_N0_364 clk__L1_N0_377 4.000000
R377_162 clk__L1_N0_366 clk__L1_N0_378 0.152000
R378_162 clk__L1_N0_366 clk__L1_N0_379 4.000000
R379_162 clk__L1_N0_367 iDFF_18_q_reg:CP 4.000000
R380_162 clk__L1_N0_368 clk__L1_N0_381 4.000000
R381_162 clk__L1_N0_370 clk__L1_N0_382 0.456000
R382_162 clk__L1_N0_371 oDFF_16_q_reg:CP 4.000000
R383_162 clk__L1_N0_373 clk__L1_N0_384 4.000000
R384_162 clk__L1_N0_374 clk__L1_N0_385 4.000000
R385_162 clk__L1_N0_375 iDFF_13_q_reg:CP 4.000000
R386_162 clk__L1_N0_376 clk__L1_N0_387 4.000000
R387_162 clk__L1_N0_377 clk_r_REG0_S2:CP 4.000000
R388_162 clk__L1_N0_378 clk__L1_N0_389 4.712000
R389_162 clk__L1_N0_378 clk__L1_N0_390 4.000000
R390_162 clk__L1_N0_379 clk__L1_N0_391 2.432000
R391_162 clk__L1_N0_381 clk__L1_N0_392 0.608000
R392_162 clk__L1_N0_382 clk__L1_N0_393 0.608000
R393_162 clk__L1_N0_382 clk__L1_N0_394 4.000000
R394_162 clk__L1_N0_384 clk__L1_N0_395 2.128000
R395_162 clk__L1_N0_385 clk_r_REG23_S2:CP 4.000000
R396_162 clk__L1_N0_387 clk__L1_N0_397 1.520000
R397_162 clk__L1_N0_389 clk__L1_N0_398 2.736000
R398_162 clk__L1_N0_389 clk__L1_N0_399 4.000000
R399_162 clk__L1_N0_389 clk__L1_N0_400 4.000000
R400_162 clk__L1_N0_390 clk_r_REG37_S2:CP 4.000000
R401_162 clk__L1_N0_391 clk__L1_N0_402 4.000000
R402_162 clk__L1_N0_392 clk__L1_N0_403 4.000000
R403_162 clk__L1_N0_393 clk__L1_N0_404 4.000000
R404_162 clk__L1_N0_394 clk_r_REG35_S2:CP 4.000000
R405_162 clk__L1_N0_395 clk__L1_N0_406 0.760000
R406_162 clk__L1_N0_395 clk__L1_N0_407 4.000000
R407_162 clk__L1_N0_397 clk__L1_N0_408 4.000000
R408_162 clk__L1_N0_398 clk__L1_N0_409 4.000000
R409_162 clk__L1_N0_399 clk__L1_N0_410 3.952000
R410_162 clk__L1_N0_411 clk__L1_N0_399 1.672000
R411_162 clk__L1_N0_400 oDFF_18_q_reg:CP 4.000000
R412_162 clk__L1_N0_402 clk__L1_N0_413 4.000000
R413_162 clk__L1_N0_403 clk_r_REG13_S2:CP 4.000000
R414_162 clk__L1_N0_404 iDFF_16_q_reg:CP 4.000000
R415_162 clk__L1_N0_406 clk__L1_N0_416 2.584000
R416_162 clk__L1_N0_406 clk__L1_N0_417 4.000000
R417_162 clk__L1_N0_407 clk_r_REG26_S2:CP 4.000000
R418_162 clk__L1_N0_408 clk__L1_N0_419 4.000000
R419_162 clk__L1_N0_420 clk__L1_N0_409 1.520000
R420_162 clk__L1_N0_409 oDFF_22_q_reg:CP 4.000000
R421_162 clk__L1_N0_410 clk__L1_N0_422 4.000000
R422_162 clk__L1_N0_411 clk__L1_N0_423 4.000000
R423_162 clk__L1_N0_413 clk_r_REG28_S2:CP 4.000000
R424_162 clk__L1_N0_416 clk__L1_N0_425 2.432000
R425_162 clk__L1_N0_416 clk__L1_N0_426 4.000000
R426_162 clk__L1_N0_417 iDFF_9_q_reg:CP 4.000000
R427_162 clk__L1_N0_419 oDFF_9_q_reg:CP 4.000000
R428_162 clk__L1_N0_420 oDFF_6_q_reg:CP 4.000000
R429_162 clk__L1_N0_430 clk__L1_N0_422 1.368000
R430_162 clk__L1_N0_422 clk__L1_N0_431 4.408000
R431_162 clk__L1_N0_422 clk__L1_N0_432 4.000000
R432_162 clk__L1_N0_433 clk__L1_N0_423 1.520000
R433_162 clk__L1_N0_423 clk__L1_N0_434 4.000000
R434_162 clk__L1_N0_425 clk__L1_N0_435 1.672000
R435_162 clk__L1_N0_425 clk__L1_N0_436 4.000000
R436_162 clk__L1_N0_426 iDFF_12_q_reg:CP 4.000000
R437_162 clk__L1_N0_430 clk__L1_N0_438 4.000000
R438_162 clk__L1_N0_431 clk__L1_N0_439 4.000000
R439_162 clk__L1_N0_432 clk_r_REG41_S2:CP 4.000000
R440_162 clk__L1_N0_433 clk__L1_N0_441 4.000000
R441_162 clk__L1_N0_434 clk_r_REG6_S2:CP 4.000000
R442_162 clk__L1_N0_435 clk__L1_N0_443 0.912000
R443_162 clk__L1_N0_435 clk__L1_N0_444 4.000000
R444_162 clk__L1_N0_445 clk__L1_N0_436 1.672000
R445_162 clk__L1_N0_438 iDFF_40_q_reg:CP 4.000000
R446_162 clk__L1_N0_439 iDFF_22_q_reg:CP 4.000000
R447_162 clk__L1_N0_441 iDFF_35_q_reg:CP 4.000000
R448_162 clk__L1_N0_443 clk__L1_N0_449 4.000000
R449_162 clk__L1_N0_444 clk__L1_N0_450 2.280000
R450_162 clk__L1_N0_445 clk__L1_N0_451 4.000000
R451_162 clk__L1_N0_449 clk_r_REG29_S2:CP 4.000000
R452_162 clk__L1_N0_450 clk__L1_N0_453 5.624000
R453_162 clk__L1_N0_450 clk__L1_N0_454 4.000000
R454_162 clk__L1_N0_451 clk__L1_N0_455 1.064000
R455_162 clk__L1_N0_451 clk__L1_N0_456 4.000000
R456_162 clk__L1_N0_453 clk__L1_N0_457 4.000000
R457_162 clk__L1_N0_454 clk__L1_N0_458 4.000000
R458_162 clk__L1_N0_455 clk__L1_N0_459 4.000000
R459_162 clk__L1_N0_456 clk_r_REG31_S2:CP 4.000000
R460_162 clk__L1_N0_461 clk__L1_N0_457 1.368000
R461_162 clk__L1_N0_458 iDFF_10_q_reg:CP 4.000000
R462_162 clk__L1_N0_463 clk__L1_N0_459 2.280000
R463_162 clk__L1_N0_461 clk__L1_N0_464 4.000000
R464_162 clk__L1_N0_465 clk__L1_N0_463 1.520000
R465_162 clk__L1_N0_463 clk__L1_N0_466 4.000000
R466_162 clk__L1_N0_464 iDFF_36_q_reg:CP 4.000000
R467_162 clk__L1_N0_465 clk__L1_N0_468 4.000000
R468_162 clk__L1_N0_466 clk__L1_N0_469 0.608000
R469_162 clk__L1_N0_466 clk__L1_N0_470 4.000000
R470_162 clk__L1_N0_468 clk__L1_N0_471 4.000000
R471_162 clk__L1_N0_469 clk__L1_N0_472 4.000000
R472_162 clk__L1_N0_470 oDFF_12_q_reg:CP 4.000000
R473_162 clk__L1_N0_471 clk__L1_I0:Z 1.000000
R474_162 clk__L1_N0_472 iDFF_14_q_reg:CP 4.000000
R475_162 clk__L1_I0:Z clk__L1_N0_476 1.000000
R476_162 clk__L1_N0_476 clk__L1_N0_477 1.368000
R477_162 clk__L1_N0_477 clk__L1_N0_478 4.000000
R478_162 clk__L1_N0_477 oDFF_10_q_reg:CP 4.000000
R479_162 clk__L1_N0_478 clk__L1_N0_480 0.304000
R480_162 clk__L1_N0_480 clk__L1_N0_481 1.976000
R481_162 clk__L1_N0_480 clk__L1_N0_482 4.000000
R482_162 clk__L1_N0_481 clk__L1_N0_483 4.000000
R483_162 clk__L1_N0_481 clk__L1_N0_484 4.000000
R484_162 clk__L1_N0_482 clk__L1_N0_485 2.280000
R485_162 clk__L1_N0_486 clk__L1_N0_483 1.672000
R486_162 clk__L1_N0_484 oDFF_14_q_reg:CP 4.000000
R487_162 clk__L1_N0_485 clk__L1_N0_488 1.672000
R488_162 clk__L1_N0_485 clk__L1_N0_489 4.000000
R489_162 clk__L1_N0_486 clk__L1_N0_490 4.000000
R490_162 clk__L1_N0_488 clk__L1_N0_491 4.000000
R491_162 clk__L1_N0_489 clk__L1_N0_492 1.064000
R492_162 clk__L1_N0_490 clk__L1_N0_493 1.520000
R493_162 clk__L1_N0_491 clk__L1_N0_494 4.560000
R494_162 clk__L1_N0_491 clk__L1_N0_495 4.000000
R495_162 clk__L1_N0_492 clk__L1_N0_496 4.000000
R496_162 clk__L1_N0_493 clk__L1_N0_497 2.280000
R497_162 clk__L1_N0_493 clk__L1_N0_498 4.000000
R498_162 clk__L1_N0_494 clk__L1_N0_499 4.000000
R499_162 clk__L1_N0_495 clk_r_REG19_S2:CP 4.000000
R500_162 clk__L1_N0_496 clk_r_REG33_S2:CP 4.000000
R501_162 clk__L1_N0_497 clk__L1_N0_502 3.496000
R502_162 clk__L1_N0_497 clk__L1_N0_503 4.000000
R503_162 clk__L1_N0_497 clk__L1_N0_504 4.000000
R504_162 clk__L1_N0_498 iDFF_11_q_reg:CP 4.000000
R505_162 clk__L1_N0_499 clk_r_REG20_S2:CP 4.000000
R506_162 clk__L1_N0_502 clk__L1_N0_507 4.000000
R507_162 clk__L1_N0_503 clk__L1_N0_508 1.672000
R508_162 clk__L1_N0_504 clk_r_REG30_S2:CP 4.000000
R509_162 clk__L1_N0_507 oDFF_11_q_reg:CP 4.000000
R510_162 clk__L1_N0_508 clk__L1_N0_511 4.000000
R511_162 clk__L1_N0_511 clk__L1_N0_512 0.608000
R512_162 clk__L1_N0_512 clk__L1_N0_513 4.000000
R513_162 clk__L1_N0_512 clk__L1_N0_514 4.000000
R514_162 clk__L1_N0_513 clk__L1_N0_515 2.280000
R515_162 clk__L1_N0_514 iDFF_15_q_reg:CP 4.000000
R516_162 clk__L1_N0_515 clk__L1_N0_517 1.672000
R517_162 clk__L1_N0_515 clk__L1_N0_518 4.000000
R518_162 clk__L1_N0_517 clk__L1_N0_519 2.280000
R519_162 clk__L1_N0_517 clk__L1_N0_520 4.000000
R520_162 clk__L1_N0_518 clk__L1_N0_521 4.000000
R521_162 clk__L1_N0_519 clk__L1_N0_522 3.952000
R522_162 clk__L1_N0_519 clk__L1_N0_523 4.000000
R523_162 clk__L1_N0_520 clk__L1_N0_524 2.888000
R524_162 clk__L1_N0_521 clk_r_REG34_S2:CP 4.000000
R525_162 clk__L1_N0_522 clk__L1_N0_526 1.672000
R526_162 clk__L1_N0_522 clk__L1_N0_527 4.000000
R527_162 clk__L1_N0_523 clk__L1_N0_528 4.000000
R528_162 clk__L1_N0_524 clk__L1_N0_529 1.672000
R529_162 clk__L1_N0_524 clk__L1_N0_530 4.000000
R530_162 clk__L1_N0_526 clk__L1_N0_531 4.000000
R531_162 clk__L1_N0_527 clk__L1_N0_532 2.432000
R532_162 clk__L1_N0_528 iDFF_2_q_reg:CP 4.000000
R533_162 clk__L1_N0_529 clk__L1_N0_534 1.368000
R534_162 clk__L1_N0_529 clk__L1_N0_535 4.000000
R535_162 clk__L1_N0_530 clk_r_REG9_S2:CP 4.000000
R536_162 clk__L1_N0_537 clk__L1_N0_531 0.608000
R537_162 clk__L1_N0_532 clk__L1_N0_538 0.456000
R538_162 clk__L1_N0_532 clk__L1_N0_539 4.000000
R539_162 clk__L1_N0_534 clk__L1_N0_540 0.152000
R540_162 clk__L1_N0_534 clk__L1_N0_541 4.000000
R541_162 clk__L1_N0_535 clk__L1_N0_542 2.280000
R542_162 clk__L1_N0_537 clk__L1_N0_543 4.000000
R543_162 clk__L1_N0_538 clk__L1_N0_544 2.432000
R544_162 clk__L1_N0_538 clk__L1_N0_545 4.000000
R545_162 clk__L1_N0_546 clk__L1_N0_539 2.280000
R546_162 clk__L1_N0_547 clk__L1_N0_540 0.304000
R547_162 clk__L1_N0_548 clk__L1_N0_541 3.952000
R548_162 clk__L1_N0_542 clk__L1_N0_549 4.000000
R549_162 clk__L1_N0_543 iDFF_6_q_reg:CP 4.000000
R550_162 clk__L1_N0_544 clk__L1_N0_551 0.152000
R551_162 clk__L1_N0_545 clk_r_REG5_S2:CP 4.000000
R552_162 clk__L1_N0_546 clk__L1_N0_553 4.000000
R553_162 clk__L1_N0_547 clk__L1_N0_554 4.000000
R554_162 clk__L1_N0_548 clk__L1_N0_555 4.000000
R555_162 clk__L1_N0_549 clk__L1_N0_556 4.000000
R556_162 clk__L1_N0_551 clk__L1_N0_557 0.304000
R557_162 clk__L1_N0_558 clk__L1_N0_553 0.304000
R558_162 clk__L1_N0_554 oDFF_2_q_reg:CP 4.000000
R559_162 clk__L1_N0_555 clk__L1_N0_560 0.304000
R560_162 clk__L1_N0_556 iDFF_3_q_reg:CP 4.000000
R561_162 clk__L1_N0_557 clk__L1_N0_562 4.000000
R562_162 clk__L1_N0_557 clk__L1_N0_563 4.000000
R563_162 clk__L1_N0_558 clk__L1_N0_564 4.000000
R564_162 clk__L1_N0_560 clk__L1_N0_565 4.000000
R565_162 clk__L1_N0_566 clk__L1_N0_562 2.432000
R566_162 clk__L1_N0_563 oDFF_7_q_reg:CP 4.000000
R567_162 clk__L1_N0_564 clk_r_REG10_S2:CP 4.000000
R568_162 clk__L1_N0_565 oDFF_15_q_reg:CP 4.000000
R569_162 clk__L1_N0_570 clk__L1_N0_566 1.520000
R570_162 clk__L1_N0_566 clk__L1_N0_571 4.000000
R571_162 clk__L1_N0_570 clk__L1_N0_572 4.000000
R572_162 clk__L1_N0_571 clk__L1_N0_573 1.368000
R573_162 clk__L1_N0_572 clk__L1_N0_574 4.000000
R574_162 clk__L1_N0_573 clk__L1_N0_575 4.000000
R575_162 clk__L1_N0_574 oDFF_3_q_reg:CP 4.000000
R576_162 clk__L1_N0_575 iDFF_7_q_reg:CP 4.000000

C1_132 oDFF_18_q_reg:Q 0 0.000045PF
C2_132 Qout_PNN741_7 0 0.000121PF
C3_132 Qout_PNN741_6 0 0.003880PF
C4_132 Qout_PNN741_5 0 0.003880PF
C5_132 Qout_PNN741_4 0 0.000111PF
C6_132 Qout_PNN741_3 0 0.000145PF
C7_132 Qout_PNN741_2 0 0.000086PF
C8_132 Qout_PNN741 0 0.000042PF
R1_132 Qout_PNN741 Qout_PNN741_2 4.000000
R2_132 Qout_PNN741_3 Qout_PNN741_2 0.152000
R3_132 Qout_PNN741_3 Qout_PNN741_4 0.912000
R4_132 Qout_PNN741_4 Qout_PNN741_5 4.000000
R5_132 Qout_PNN741_6 Qout_PNN741_5 33.135999
R6_132 Qout_PNN741_6 Qout_PNN741_7 4.000000
R7_132 Qout_PNN741_7 oDFF_18_q_reg:Q 4.000000

C1_120 oDFF_6_q_reg:Q 0 0.000045PF
C2_120 Qout_PNN729_7 0 0.000044PF
C3_120 Qout_PNN729_6 0 0.000044PF
C4_120 Qout_PNN729_5 0 0.003585PF
C5_120 Qout_PNN729_4 0 0.003585PF
C6_120 Qout_PNN729_3 0 0.000067PF
C7_120 Qout_PNN729_2 0 0.000067PF
C8_120 Qout_PNN729 0 0.000042PF
R1_120 Qout_PNN729 Qout_PNN729_2 4.000000
R2_120 Qout_PNN729_3 Qout_PNN729_2 0.608000
R3_120 Qout_PNN729_3 Qout_PNN729_4 4.000000
R4_120 Qout_PNN729_5 Qout_PNN729_4 30.551999
R5_120 Qout_PNN729_5 Qout_PNN729_6 4.000000
R6_120 Qout_PNN729_7 Qout_PNN729_6 0.304000
R7_120 Qout_PNN729_7 oDFF_6_q_reg:Q 4.000000

C1_74 PNN69 0 0.000042PF
C2_74 PNN69_7 0 0.000104PF
C3_74 PNN69_6 0 0.000104PF
C4_74 PNN69_5 0 0.005036PF
C5_74 PNN69_4 0 0.005036PF
C6_74 PNN69_3 0 0.000050PF
C7_74 PNN69_2 0 0.000034PF
C8_74 iDFF_18_q_reg:D 0 0.000045PF
R1_74 iDFF_18_q_reg:D PNN69_2 4.000000
R2_74 PNN69_2 PNN69_3 0.152000
R3_74 PNN69_3 PNN69_4 4.000000
R4_74 PNN69_4 PNN69_5 40.735999
R5_74 PNN69_5 PNN69_6 4.000000
R6_74 PNN69_7 PNN69_6 0.304000
R7_74 PNN69_7 PNN69 4.000000

C1_135 oDFF_21_q_reg:Q 0 0.000045PF
C2_135 Qout_PNN744_7 0 0.000044PF
C3_135 Qout_PNN744_6 0 0.000044PF
C4_135 Qout_PNN744_5 0 0.002436PF
C5_135 Qout_PNN744_4 0 0.002436PF
C6_135 Qout_PNN744_3 0 0.000056PF
C7_135 Qout_PNN744_2 0 0.000056PF
C8_135 Qout_PNN744 0 0.000042PF
R1_135 Qout_PNN744 Qout_PNN744_2 4.000000
R2_135 Qout_PNN744_3 Qout_PNN744_2 0.456000
R3_135 Qout_PNN744_3 Qout_PNN744_4 4.000000
R4_135 Qout_PNN744_5 Qout_PNN744_4 30.551999
R5_135 Qout_PNN744_5 Qout_PNN744_6 4.000000
R6_135 Qout_PNN744_7 Qout_PNN744_6 0.304000
R7_135 Qout_PNN744_7 oDFF_21_q_reg:Q 4.000000

C1_138 oDFF_24_q_reg:Q 0 0.000045PF
C2_138 Qout_PNN747_7 0 0.000044PF
C3_138 Qout_PNN747_6 0 0.000044PF
C4_138 Qout_PNN747_5 0 0.002511PF
C5_138 Qout_PNN747_4 0 0.002511PF
C6_138 Qout_PNN747_3 0 0.000044PF
C7_138 Qout_PNN747_2 0 0.000044PF
C8_138 Qout_PNN747 0 0.000042PF
R1_138 Qout_PNN747 Qout_PNN747_2 4.000000
R2_138 Qout_PNN747_2 Qout_PNN747_3 0.304000
R3_138 Qout_PNN747_3 Qout_PNN747_4 4.000000
R4_138 Qout_PNN747_5 Qout_PNN747_4 30.551999
R5_138 Qout_PNN747_5 Qout_PNN747_6 4.000000
R6_138 Qout_PNN747_7 Qout_PNN747_6 0.304000
R7_138 Qout_PNN747_7 oDFF_24_q_reg:Q 4.000000

C1_54 PNN132 0 0.000084PF
C2_54 PNN132_17 0 0.000216PF
C3_54 PNN132_16 0 0.000093PF
C4_54 PNN132_15 0 0.003075PF
C5_54 PNN132_14 0 0.003075PF
C6_54 PNN132_13 0 0.000052PF
C7_54 PNN132_12 0 0.000036PF
C8_54 PNN132_11 0 0.000713PF
C9_54 PNN132_10 0 0.000713PF
C10_54 PNN132_9 0 0.000054PF
C11_54 PNN132_8 0 0.000071PF
C12_54 PNN132_7 0 0.001263PF
C13_54 PNN132_6 0 0.001263PF
C14_54 PNN132_5 0 0.000231PF
C15_54 PNN132_4 0 0.000231PF
C16_54 PNN132_3 0 0.000072PF
C17_54 PNN132_2 0 0.000072PF
C18_54 iDFF_36_q_reg:D 0 0.000045PF
R1_54 iDFF_36_q_reg:D PNN132_2 4.000000
R2_54 PNN132_3 PNN132_2 0.608000
R3_54 PNN132_3 PNN132_4 4.000000
R4_54 PNN132_4 PNN132_5 1.064000
R5_54 PNN132_5 PNN132_6 4.000000
R6_54 PNN132_7 PNN132_6 8.968000
R7_54 PNN132_7 PNN132_8 4.000000
R8_54 PNN132_8 PNN132_9 0.152000
R9_54 PNN132_9 PNN132_10 4.000000
R10_54 PNN132_11 PNN132_10 3.648000
R11_54 PNN132_11 PNN132_12 4.000000
R12_54 PNN132_13 PNN132_12 0.152000
R13_54 PNN132_13 PNN132_14 4.000000
R14_54 PNN132_15 PNN132_14 31.007999
R15_54 PNN132_15 PNN132_16 4.000000
R16_54 PNN132_17 PNN132_16 0.528000
R17_54 PNN132_17 PNN132 4.000000

C1_63 PNN29 0 0.000042PF
C2_63 PNN29_11 0 0.000121PF
C3_63 PNN29_10 0 0.001593PF
C4_63 PNN29_9 0 0.001593PF
C5_63 PNN29_8 0 0.000121PF
C6_63 PNN29_7 0 0.001843PF
C7_63 PNN29_6 0 0.001877PF
C8_63 PNN29_5 0 0.000255PF
C9_63 PNN29_4 0 0.000221PF
C10_63 PNN29_3 0 0.000064PF
C11_63 PNN29_2 0 0.000064PF
C12_63 iDFF_8_q_reg:D 0 0.000045PF
R1_63 iDFF_8_q_reg:D PNN29_2 4.000000
R2_63 PNN29_3 PNN29_2 0.304000
R3_63 PNN29_3 PNN29_4 4.000000
R4_63 PNN29_5 PNN29_4 2.736000
R5_63 PNN29_5 PNN29_6 0.152000
R6_63 PNN29_7 PNN29_6 22.951999
R7_63 PNN29_7 PNN29_8 4.000000
R8_63 PNN29_8 PNN29_9 4.000000
R9_63 PNN29_10 PNN29_9 4.136000
R10_63 PNN29_10 PNN29_11 4.000000
R11_63 PNN29_11 PNN29 4.000000

C1_115 oDFF_1_q_reg:Q 0 0.000045PF
C2_115 Qout_PNN724_10 0 0.000033PF
C3_115 Qout_PNN724_9 0 0.000049PF
C4_115 Qout_PNN724_8 0 0.000121PF
C5_115 Qout_PNN724_7 0 0.000033PF
C6_115 Qout_PNN724_6 0 0.000049PF
C7_115 Qout_PNN724_5 0 0.003403PF
C8_115 Qout_PNN724_4 0 0.003403PF
C9_115 Qout_PNN724_3 0 0.000044PF
C10_115 Qout_PNN724_2 0 0.000044PF
C11_115 Qout_PNN724 0 0.000042PF
R1_115 Qout_PNN724 Qout_PNN724_2 4.000000
R2_115 Qout_PNN724_2 Qout_PNN724_3 0.304000
R3_115 Qout_PNN724_3 Qout_PNN724_4 4.000000
R4_115 Qout_PNN724_4 Qout_PNN724_5 17.688000
R5_115 Qout_PNN724_5 Qout_PNN724_6 4.000000
R6_115 Qout_PNN724_7 Qout_PNN724_6 0.152000
R7_115 Qout_PNN724_7 Qout_PNN724_8 4.000000
R8_115 Qout_PNN724_8 Qout_PNN724_9 4.000000
R9_115 Qout_PNN724_10 Qout_PNN724_9 0.152000
R10_115 Qout_PNN724_10 oDFF_1_q_reg:Q 4.000000

C1_51 PNN13 0 0.002317PF
C2_51 PNN13_6 0 0.002338PF
C3_51 PNN13_5 0 0.000121PF
C4_51 PNN13_4 0 0.000178PF
C5_51 PNN13_3 0 0.000178PF
C6_51 PNN13_2 0 0.000121PF
C7_51 iDFF_4_q_reg:D 0 0.000045PF
R1_51 iDFF_4_q_reg:D PNN13_2 4.000000
R2_51 PNN13_2 PNN13_3 4.000000
R3_51 PNN13_4 PNN13_3 1.368000
R4_51 PNN13_4 PNN13_5 4.000000
R5_51 PNN13_5 PNN13_6 4.000000
R6_51 PNN13 PNN13_6 16.808000

C1_118 oDFF_4_q_reg:Q 0 0.000045PF
C2_118 Qout_PNN727_8 0 0.000121PF
C3_118 Qout_PNN727_7 0 0.001861PF
C4_118 Qout_PNN727_6 0 0.001861PF
C5_118 Qout_PNN727_5 0 0.000121PF
C6_118 Qout_PNN727_4 0 0.000598PF
C7_118 Qout_PNN727_3 0 0.000598PF
C8_118 Qout_PNN727_2 0 0.000121PF
C9_118 Qout_PNN727 0 0.000042PF
R1_118 Qout_PNN727 Qout_PNN727_2 4.000000
R2_118 Qout_PNN727_2 Qout_PNN727_3 4.000000
R3_118 Qout_PNN727_3 Qout_PNN727_4 4.224000
R4_118 Qout_PNN727_4 Qout_PNN727_5 4.000000
R5_118 Qout_PNN727_5 Qout_PNN727_6 4.000000
R6_118 Qout_PNN727_6 Qout_PNN727_7 23.255999
R7_118 Qout_PNN727_7 Qout_PNN727_8 4.000000
R8_118 Qout_PNN727_8 oDFF_4_q_reg:Q 4.000000

C1_121 oDFF_7_q_reg:Q 0 0.000045PF
C2_121 Qout_PNN730_11 0 0.000121PF
C3_121 Qout_PNN730_10 0 0.000513PF
C4_121 Qout_PNN730_9 0 0.000548PF
C5_121 Qout_PNN730_8 0 0.001298PF
C6_121 Qout_PNN730_7 0 0.001263PF
C7_121 Qout_PNN730_6 0 0.000121PF
C8_121 Qout_PNN730_5 0 0.000742PF
C9_121 Qout_PNN730_4 0 0.000742PF
C10_121 Qout_PNN730_3 0 0.000049PF
C11_121 Qout_PNN730_2 0 0.000032PF
C12_121 Qout_PNN730 0 0.000042PF
R1_121 Qout_PNN730 Qout_PNN730_2 4.000000
R2_121 Qout_PNN730_3 Qout_PNN730_2 0.152000
R3_121 Qout_PNN730_3 Qout_PNN730_4 4.000000
R4_121 Qout_PNN730_5 Qout_PNN730_4 5.280000
R5_121 Qout_PNN730_5 Qout_PNN730_6 4.000000
R6_121 Qout_PNN730_6 Qout_PNN730_7 4.000000
R7_121 Qout_PNN730_8 Qout_PNN730_7 15.200000
R8_121 Qout_PNN730_8 Qout_PNN730_9 0.152000
R9_121 Qout_PNN730_10 Qout_PNN730_9 6.232000
R10_121 Qout_PNN730_10 Qout_PNN730_11 4.000000
R11_121 Qout_PNN730_11 oDFF_7_q_reg:Q 4.000000

C1_61 PNN21 0 0.000042PF
C2_61 PNN21_9 0 0.000121PF
C3_61 PNN21_8 0 0.000782PF
C4_61 PNN21_7 0 0.000782PF
C5_61 PNN21_6 0 0.000121PF
C6_61 PNN21_5 0 0.002050PF
C7_61 PNN21_4 0 0.002050PF
C8_61 PNN21_3 0 0.000121PF
C9_61 PNN21_2 0 0.000362PF
C10_61 iDFF_6_q_reg:D 0 0.000340PF
R1_61 iDFF_6_q_reg:D PNN21_2 3.648000
R2_61 PNN21_2 PNN21_3 4.000000
R3_61 PNN21_3 PNN21_4 4.000000
R4_61 PNN21_4 PNN21_5 25.535999
R5_61 PNN21_5 PNN21_6 4.000000
R6_61 PNN21_6 PNN21_7 4.000000
R7_61 PNN21_7 PNN21_8 5.368000
R8_61 PNN21_8 PNN21_9 4.000000
R9_61 PNN21_9 PNN21 4.000000

C1_55 PNN133 0 0.002996PF
C2_55 PNN133_6 0 0.003017PF
C3_55 PNN133_5 0 0.000121PF
C4_55 PNN133_4 0 0.001621PF
C5_55 PNN133_3 0 0.001621PF
C6_55 PNN133_2 0 0.000121PF
C7_55 iDFF_37_q_reg:D 0 0.000045PF
R1_55 iDFF_37_q_reg:D PNN133_2 4.000000
R2_55 PNN133_2 PNN133_3 4.000000
R3_55 PNN133_3 PNN133_4 6.080000
R4_55 PNN133_4 PNN133_5 4.000000
R5_55 PNN133_5 PNN133_6 4.000000
R6_55 PNN133_6 PNN133 21.736000

C1_59 PNN137 0 0.007787PF
C2_59 PNN137_6 0 0.007808PF
C3_59 PNN137_5 0 0.000071PF
C4_59 PNN137_4 0 0.000055PF
C5_59 PNN137_3 0 0.000121PF
C6_59 PNN137_2 0 0.000121PF
C7_59 iDFF_41_q_reg:D 0 0.000045PF
R1_59 iDFF_41_q_reg:D PNN137_2 4.000000
R2_59 PNN137_2 PNN137_3 4.000000
R3_59 PNN137_3 PNN137_4 4.000000
R4_59 PNN137_5 PNN137_4 0.152000
R5_59 PNN137_5 PNN137_6 4.000000
R6_59 PNN137_6 PNN137 24.904000

C1_136 oDFF_22_q_reg:Q 0 0.000045PF
C2_136 Qout_PNN745_9 0 0.000045PF
C3_136 Qout_PNN745_8 0 0.000045PF
C4_136 Qout_PNN745_7 0 0.000121PF
C5_136 Qout_PNN745_6 0 0.000121PF
C6_136 Qout_PNN745_5 0 0.006845PF
C7_136 Qout_PNN745_4 0 0.006845PF
C8_136 Qout_PNN745_3 0 0.000077PF
C9_136 Qout_PNN745_2 0 0.000077PF
C10_136 Qout_PNN745 0 0.000042PF
R1_136 Qout_PNN745 Qout_PNN745_2 4.000000
R2_136 Qout_PNN745_2 Qout_PNN745_3 0.456000
R3_136 Qout_PNN745_3 Qout_PNN745_4 4.000000
R4_136 Qout_PNN745_5 Qout_PNN745_4 17.776000
R5_136 Qout_PNN745_5 Qout_PNN745_6 4.000000
R6_136 Qout_PNN745_6 Qout_PNN745_7 4.000000
R7_136 Qout_PNN745_7 Qout_PNN745_8 4.000000
R8_136 Qout_PNN745_9 Qout_PNN745_8 0.304000
R9_136 Qout_PNN745_9 oDFF_22_q_reg:Q 4.000000

C1_57 PNN135 0 0.000042PF
C2_57 PNN135_19 0 0.000121PF
C3_57 PNN135_18 0 0.000563PF
C4_57 PNN135_17 0 0.000563PF
C5_57 PNN135_16 0 0.000121PF
C6_57 PNN135_15 0 0.002903PF
C7_57 PNN135_14 0 0.002903PF
C8_57 PNN135_13 0 0.000121PF
C9_57 PNN135_12 0 0.000540PF
C10_57 PNN135_11 0 0.000540PF
C11_57 PNN135_10 0 0.000121PF
C12_57 PNN135_9 0 0.000464PF
C13_57 PNN135_8 0 0.000464PF
C14_57 PNN135_7 0 0.000050PF
C15_57 PNN135_6 0 0.000050PF
C16_57 PNN135_5 0 0.000801PF
C17_57 PNN135_4 0 0.000801PF
C18_57 PNN135_3 0 0.000056PF
C19_57 PNN135_2 0 0.000056PF
C20_57 iDFF_39_q_reg:D 0 0.000045PF
R1_57 iDFF_39_q_reg:D PNN135_2 4.000000
R2_57 PNN135_3 PNN135_2 0.304000
R3_57 PNN135_3 PNN135_4 4.000000
R4_57 PNN135_5 PNN135_4 4.408000
R5_57 PNN135_5 PNN135_6 4.000000
R6_57 PNN135_6 PNN135_7 0.304000
R7_57 PNN135_7 PNN135_8 4.000000
R8_57 PNN135_9 PNN135_8 1.216000
R9_57 PNN135_9 PNN135_10 4.000000
R10_57 PNN135_10 PNN135_11 4.000000
R11_57 PNN135_12 PNN135_11 3.960000
R12_57 PNN135_12 PNN135_13 4.000000
R13_57 PNN135_13 PNN135_14 4.000000
R14_57 PNN135_15 PNN135_14 25.687999
R15_57 PNN135_15 PNN135_16 4.000000
R16_57 PNN135_16 PNN135_17 4.000000
R17_57 PNN135_18 PNN135_17 4.136000
R18_57 PNN135_18 PNN135_19 4.000000
R19_57 PNN135_19 PNN135 4.000000

C1_58 PNN136 0 0.002853PF
C2_58 PNN136_6 0 0.002874PF
C3_58 PNN136_5 0 0.000049PF
C4_58 PNN136_4 0 0.000032PF
C5_58 PNN136_3 0 0.000121PF
C6_58 PNN136_2 0 0.000121PF
C7_58 iDFF_40_q_reg:D 0 0.000045PF
R1_58 iDFF_40_q_reg:D PNN136_2 4.000000
R2_58 PNN136_2 PNN136_3 4.000000
R3_58 PNN136_3 PNN136_4 4.000000
R4_58 PNN136_5 PNN136_4 0.152000
R5_58 PNN136_5 PNN136_6 4.000000
R6_58 PNN136_6 PNN136 21.032000

C1_47 PNN117 0 0.000042PF
C2_47 PNN117_8 0 0.000121PF
C3_47 PNN117_7 0 0.000622PF
C4_47 PNN117_6 0 0.000622PF
C5_47 PNN117_5 0 0.000121PF
C6_47 PNN117_4 0 0.001896PF
C7_47 PNN117_3 0 0.001896PF
C8_47 PNN117_2 0 0.000121PF
C9_47 iDFF_30_q_reg:D 0 0.000045PF
R1_47 iDFF_30_q_reg:D PNN117_2 4.000000
R2_47 PNN117_2 PNN117_3 4.000000
R3_47 PNN117_4 PNN117_3 22.799999
R4_47 PNN117_4 PNN117_5 4.000000
R5_47 PNN117_5 PNN117_6 4.000000
R6_47 PNN117_7 PNN117_6 4.400000
R7_47 PNN117_7 PNN117_8 4.000000
R8_47 PNN117_8 PNN117 4.000000

C1_43 PNN101 0 0.000042PF
C2_43 PNN101_11 0 0.000121PF
C3_43 PNN101_10 0 0.001717PF
C4_43 PNN101_9 0 0.001717PF
C5_43 PNN101_8 0 0.000121PF
C6_43 PNN101_7 0 0.001114PF
C7_43 PNN101_6 0 0.001204PF
C8_43 PNN101_5 0 0.001216PF
C9_43 PNN101_4 0 0.001126PF
C10_43 PNN101_3 0 0.000067PF
C11_43 PNN101_2 0 0.000067PF
C12_43 iDFF_26_q_reg:D 0 0.000045PF
R1_43 iDFF_26_q_reg:D PNN101_2 4.000000
R2_43 PNN101_3 PNN101_2 0.456000
R3_43 PNN101_3 PNN101_4 4.000000
R4_43 PNN101_5 PNN101_4 11.400000
R5_43 PNN101_5 PNN101_6 0.304000
R6_43 PNN101_7 PNN101_6 13.832000
R7_43 PNN101_7 PNN101_8 4.000000
R8_43 PNN101_8 PNN101_9 4.000000
R9_43 PNN101_10 PNN101_9 4.400000
R10_43 PNN101_10 PNN101_11 4.000000
R11_43 PNN101_11 PNN101 4.000000

C1_140 oDFF_26_q_reg:Q 0 0.000045PF
C2_140 Qout_PNN749_10 0 0.000045PF
C3_140 Qout_PNN749_9 0 0.000045PF
C4_140 Qout_PNN749_8 0 0.000872PF
C5_140 Qout_PNN749_7 0 0.000872PF
C6_140 Qout_PNN749_6 0 0.000121PF
C7_140 Qout_PNN749_5 0 0.002755PF
C8_140 Qout_PNN749_4 0 0.002755PF
C9_140 Qout_PNN749_3 0 0.000044PF
C10_140 Qout_PNN749_2 0 0.000044PF
C11_140 Qout_PNN749 0 0.000042PF
R1_140 Qout_PNN749 Qout_PNN749_2 4.000000
R2_140 Qout_PNN749_2 Qout_PNN749_3 0.304000
R3_140 Qout_PNN749_3 Qout_PNN749_4 4.000000
R4_140 Qout_PNN749_4 Qout_PNN749_5 12.496000
R5_140 Qout_PNN749_5 Qout_PNN749_6 4.000000
R6_140 Qout_PNN749_6 Qout_PNN749_7 4.000000
R7_140 Qout_PNN749_7 Qout_PNN749_8 8.968000
R8_140 Qout_PNN749_8 Qout_PNN749_9 4.000000
R9_140 Qout_PNN749_10 Qout_PNN749_9 0.304000
R10_140 Qout_PNN749_10 oDFF_26_q_reg:Q 4.000000



XFE_OFCC1_n168 FE_OFCC1_n168:Z FE_OFCC1_n168:A gnd gnds vdd vdds HS65_GS_BFX18
XFE_OFCC0_c0_n49 FE_OFCC0_c0_n49:Z FE_OFCC0_c0_n49:A gnd gnds vdd vdds HS65_GS_BFX18
Xclk__L1_I0 clk__L1_I0:Z clk__L1_I0:A gnd gnds vdd vdds HS65_GS_BFX284
XiDFF_1_q_reg iDFF_1_q_reg:Q iDFF_1_q_reg:D iDFF_1_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_2_q_reg iDFF_2_q_reg:Q iDFF_2_q_reg:D iDFF_2_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_3_q_reg iDFF_3_q_reg:Q iDFF_3_q_reg:D iDFF_3_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_4_q_reg iDFF_4_q_reg:Q iDFF_4_q_reg:D iDFF_4_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9_21
XiDFF_6_q_reg iDFF_6_q_reg:Q iDFF_6_q_reg:D iDFF_6_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_7_q_reg iDFF_7_q_reg:Q iDFF_7_q_reg:D iDFF_7_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_8_q_reg iDFF_8_q_reg:Q iDFF_8_q_reg:D iDFF_8_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_9_q_reg iDFF_9_q_reg:Q iDFF_9_q_reg:D iDFF_9_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_10_q_reg iDFF_10_q_reg:Q iDFF_10_q_reg:D iDFF_10_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_11_q_reg iDFF_11_q_reg:Q iDFF_11_q_reg:D iDFF_11_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_12_q_reg iDFF_12_q_reg:Q iDFF_12_q_reg:D iDFF_12_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_13_q_reg iDFF_13_q_reg:Q iDFF_13_q_reg:D iDFF_13_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_14_q_reg iDFF_14_q_reg:Q iDFF_14_q_reg:D iDFF_14_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_15_q_reg iDFF_15_q_reg:Q iDFF_15_q_reg:D iDFF_15_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_16_q_reg iDFF_16_q_reg:Q iDFF_16_q_reg:D iDFF_16_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_17_q_reg iDFF_17_q_reg:Q iDFF_17_q_reg:D iDFF_17_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_18_q_reg iDFF_18_q_reg:Q iDFF_18_q_reg:D iDFF_18_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_19_q_reg iDFF_19_q_reg:Q iDFF_19_q_reg:D iDFF_19_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_20_q_reg iDFF_20_q_reg:Q iDFF_20_q_reg:D iDFF_20_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_21_q_reg iDFF_21_q_reg:Q iDFF_21_q_reg:D iDFF_21_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_22_q_reg iDFF_22_q_reg:Q iDFF_22_q_reg:D iDFF_22_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_23_q_reg iDFF_23_q_reg:Q iDFF_23_q_reg:D iDFF_23_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_24_q_reg iDFF_24_q_reg:Q iDFF_24_q_reg:D iDFF_24_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_25_q_reg iDFF_25_q_reg:Q iDFF_25_q_reg:D iDFF_25_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_26_q_reg iDFF_26_q_reg:Q iDFF_26_q_reg:D iDFF_26_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_27_q_reg iDFF_27_q_reg:Q iDFF_27_q_reg:D iDFF_27_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_28_q_reg iDFF_28_q_reg:Q iDFF_28_q_reg:D iDFF_28_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_29_q_reg iDFF_29_q_reg:Q iDFF_29_q_reg:D iDFF_29_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_30_q_reg iDFF_30_q_reg:Q iDFF_30_q_reg:D iDFF_30_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_31_q_reg iDFF_31_q_reg:Q iDFF_31_q_reg:D iDFF_31_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_32_q_reg iDFF_32_q_reg:Q iDFF_32_q_reg:D iDFF_32_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_33_q_reg iDFF_33_q_reg:Q iDFF_33_q_reg:D iDFF_33_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_34_q_reg iDFF_34_q_reg:Q iDFF_34_q_reg:D iDFF_34_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_35_q_reg iDFF_35_q_reg:Q iDFF_35_q_reg:D iDFF_35_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_36_q_reg iDFF_36_q_reg:Q iDFF_36_q_reg:D iDFF_36_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_37_q_reg iDFF_37_q_reg:Q iDFF_37_q_reg:D iDFF_37_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_38_q_reg iDFF_38_q_reg:Q iDFF_38_q_reg:D iDFF_38_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_39_q_reg iDFF_39_q_reg:Q iDFF_39_q_reg:D iDFF_39_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_40_q_reg iDFF_40_q_reg:Q iDFF_40_q_reg:D iDFF_40_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_41_q_reg iDFF_41_q_reg:Q iDFF_41_q_reg:D iDFF_41_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_1_q_reg oDFF_1_q_reg:Q oDFF_1_q_reg:D oDFF_1_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_2_q_reg oDFF_2_q_reg:Q oDFF_2_q_reg:D oDFF_2_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_3_q_reg oDFF_3_q_reg:Q oDFF_3_q_reg:D oDFF_3_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_4_q_reg oDFF_4_q_reg:Q oDFF_4_q_reg:D oDFF_4_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_5_q_reg oDFF_5_q_reg:Q oDFF_5_q_reg:D oDFF_5_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_6_q_reg oDFF_6_q_reg:Q oDFF_6_q_reg:D oDFF_6_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_7_q_reg oDFF_7_q_reg:Q oDFF_7_q_reg:D oDFF_7_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_8_q_reg oDFF_8_q_reg:Q oDFF_8_q_reg:D oDFF_8_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_9_q_reg oDFF_9_q_reg:Q oDFF_9_q_reg:D oDFF_9_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_10_q_reg oDFF_10_q_reg:Q oDFF_10_q_reg:D oDFF_10_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_11_q_reg oDFF_11_q_reg:Q oDFF_11_q_reg:D oDFF_11_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_12_q_reg oDFF_12_q_reg:Q oDFF_12_q_reg:D oDFF_12_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_13_q_reg oDFF_13_q_reg:Q oDFF_13_q_reg:D oDFF_13_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_14_q_reg oDFF_14_q_reg:Q oDFF_14_q_reg:D oDFF_14_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_15_q_reg oDFF_15_q_reg:Q oDFF_15_q_reg:D oDFF_15_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_16_q_reg oDFF_16_q_reg:Q oDFF_16_q_reg:D oDFF_16_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_17_q_reg oDFF_17_q_reg:Q oDFF_17_q_reg:D oDFF_17_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_18_q_reg oDFF_18_q_reg:Q oDFF_18_q_reg:D oDFF_18_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_19_q_reg oDFF_19_q_reg:Q oDFF_19_q_reg:D oDFF_19_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_20_q_reg oDFF_20_q_reg:Q oDFF_20_q_reg:D oDFF_20_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_21_q_reg oDFF_21_q_reg:Q oDFF_21_q_reg:D oDFF_21_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_22_q_reg oDFF_22_q_reg:Q oDFF_22_q_reg:D oDFF_22_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_23_q_reg oDFF_23_q_reg:Q oDFF_23_q_reg:D oDFF_23_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_24_q_reg oDFF_24_q_reg:Q oDFF_24_q_reg:D oDFF_24_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_25_q_reg oDFF_25_q_reg:Q oDFF_25_q_reg:D oDFF_25_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_26_q_reg oDFF_26_q_reg:Q oDFF_26_q_reg:D oDFF_26_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_27_q_reg oDFF_27_q_reg:Q oDFF_27_q_reg:D oDFF_27_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_28_q_reg oDFF_28_q_reg:Q oDFF_28_q_reg:D oDFF_28_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_29_q_reg oDFF_29_q_reg:Q oDFF_29_q_reg:D oDFF_29_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_30_q_reg oDFF_30_q_reg:Q oDFF_30_q_reg:D oDFF_30_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_31_q_reg oDFF_31_q_reg:Q oDFF_31_q_reg:D oDFF_31_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XoDFF_32_q_reg oDFF_32_q_reg:Q oDFF_32_q_reg:D oDFF_32_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG28_S2 clk_r_REG28_S2:Q clk_r_REG28_S2:D clk_r_REG28_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG16_S2 clk_r_REG16_S2:Q clk_r_REG16_S2:D clk_r_REG16_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG25_S2 clk_r_REG25_S2:Q clk_r_REG25_S2:D clk_r_REG25_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG13_S2 clk_r_REG13_S2:Q clk_r_REG13_S2:D clk_r_REG13_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG1_S2 clk_r_REG1_S2:Q clk_r_REG1_S2:D clk_r_REG1_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG5_S2 clk_r_REG5_S2:Q clk_r_REG5_S2:D clk_r_REG5_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG6_S2 clk_r_REG6_S2:Q clk_r_REG6_S2:D clk_r_REG6_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG8_S2 clk_r_REG8_S2:Q clk_r_REG8_S2:D clk_r_REG8_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG9_S2 clk_r_REG9_S2:Q clk_r_REG9_S2:D clk_r_REG9_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG7_S2 clk_r_REG7_S2:Q clk_r_REG7_S2:D clk_r_REG7_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG10_S2 clk_r_REG10_S2:Q clk_r_REG10_S2:D clk_r_REG10_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG2_S2 clk_r_REG2_S2:Q clk_r_REG2_S2:D clk_r_REG2_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG21_S2 clk_r_REG21_S2:Q clk_r_REG21_S2:D clk_r_REG21_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG22_S2 clk_r_REG22_S2:Q clk_r_REG22_S2:D clk_r_REG22_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG3_S2 clk_r_REG3_S2:Q clk_r_REG3_S2:D clk_r_REG3_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG17_S2 clk_r_REG17_S2:Q clk_r_REG17_S2:D clk_r_REG17_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG18_S2 clk_r_REG18_S2:Q clk_r_REG18_S2:D clk_r_REG18_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG26_S2 clk_r_REG26_S2:Q clk_r_REG26_S2:D clk_r_REG26_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG29_S2 clk_r_REG29_S2:Q clk_r_REG29_S2:D clk_r_REG29_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG30_S2 clk_r_REG30_S2:Q clk_r_REG30_S2:D clk_r_REG30_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG31_S2 clk_r_REG31_S2:Q clk_r_REG31_S2:D clk_r_REG31_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG32_S2 clk_r_REG32_S2:Q clk_r_REG32_S2:D clk_r_REG32_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG33_S2 clk_r_REG33_S2:Q clk_r_REG33_S2:D clk_r_REG33_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG34_S2 clk_r_REG34_S2:Q clk_r_REG34_S2:D clk_r_REG34_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG35_S2 clk_r_REG35_S2:Q clk_r_REG35_S2:D clk_r_REG35_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG36_S2 clk_r_REG36_S2:Q clk_r_REG36_S2:D clk_r_REG36_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG37_S2 clk_r_REG37_S2:Q clk_r_REG37_S2:D clk_r_REG37_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG38_S2 clk_r_REG38_S2:Q clk_r_REG38_S2:D clk_r_REG38_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG39_S2 clk_r_REG39_S2:Q clk_r_REG39_S2:D clk_r_REG39_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG40_S2 clk_r_REG40_S2:Q clk_r_REG40_S2:D clk_r_REG40_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG41_S2 clk_r_REG41_S2:Q clk_r_REG41_S2:D clk_r_REG41_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG42_S2 clk_r_REG42_S2:Q clk_r_REG42_S2:D clk_r_REG42_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG43_S2 clk_r_REG43_S2:Q clk_r_REG43_S2:D clk_r_REG43_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG44_S2 clk_r_REG44_S2:Q clk_r_REG44_S2:D clk_r_REG44_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG45_S2 clk_r_REG45_S2:Q clk_r_REG45_S2:D clk_r_REG45_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG46_S2 clk_r_REG46_S2:Q clk_r_REG46_S2:D clk_r_REG46_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG47_S2 clk_r_REG47_S2:Q clk_r_REG47_S2:D clk_r_REG47_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG48_S2 clk_r_REG48_S2:Q clk_r_REG48_S2:D clk_r_REG48_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG49_S2 clk_r_REG49_S2:Q clk_r_REG49_S2:D clk_r_REG49_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG50_S2 clk_r_REG50_S2:Q clk_r_REG50_S2:D clk_r_REG50_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG51_S2 clk_r_REG51_S2:Q clk_r_REG51_S2:D clk_r_REG51_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG0_S2 clk_r_REG0_S2:Q clk_r_REG0_S2:D clk_r_REG0_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG12_S2 clk_r_REG12_S2:Q clk_r_REG12_S2:D clk_r_REG12_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG15_S2 clk_r_REG15_S2:Q clk_r_REG15_S2:D clk_r_REG15_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG27_S2 clk_r_REG27_S2:Q clk_r_REG27_S2:D clk_r_REG27_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG4_S2 clk_r_REG4_S2:Q clk_r_REG4_S2:D clk_r_REG4_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG11_S2 clk_r_REG11_S2:Q clk_r_REG11_S2:D clk_r_REG11_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG24_S2 clk_r_REG24_S2:Q clk_r_REG24_S2:D clk_r_REG24_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG20_S2 clk_r_REG20_S2:Q clk_r_REG20_S2:D clk_r_REG20_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG23_S2 clk_r_REG23_S2:Q clk_r_REG23_S2:D clk_r_REG23_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG19_S2 clk_r_REG19_S2:Q clk_r_REG19_S2:D clk_r_REG19_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
Xclk_r_REG14_S2 clk_r_REG14_S2:Q clk_r_REG14_S2:D clk_r_REG14_S2:CP gnd gnds vdd vdds HS65_GS_DFPQX9
XiDFF_5_q_reg iDFF_5_q_reg:QN iDFF_5_q_reg:D iDFF_5_q_reg:CP gnd gnds vdd vdds HS65_GS_DFPQNX9
XU159 U159:Z U159:C U159:B U159:A gnd gnds vdd vdds HS65_GSS_XOR3X4
XU160 U160:Z U160:C U160:B U160:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU161 U161:Z U161:B U161:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU162 U162:Z U162:C U162:B U162:A gnd gnds vdd vdds HS65_GS_NOR3X4
XU163 U163:Z U163:B U163:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU164 U164:Z U164:B U164:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU165 U165:Z U165:B U165:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU166 U166:Z U166:E U166:D U166:C U166:B U166:A gnd gnds vdd vdds HS65_GS_OAI32X5
XU167 U167:Z U167:C U167:B U167:A gnd gnds vdd vdds HS65_GS_AOI12X2
XU168 U168:Z U168:C U168:B U168:A gnd gnds vdd vdds HS65_GS_AOI12X2
XU169 U169:Z U169:E U169:D U169:C U169:B U169:A gnd gnds vdd vdds HS65_GS_AOI32X5
XU170 U170:Z U170:P U170:B U170:A gnd gnds vdd vdds HS65_GS_PAOI2X1
XU171 U171:Z U171:C U171:B U171:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU172 U172:Z U172:C U172:B U172:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU173 U173:Z U173:C U173:B U173:A gnd gnds vdd vdds HS65_GSS_XOR3X4
XU174 U174:Z U174:B U174:A gnd gnds vdd vdds HS65_GSS_XNOR2X6
XU175 U175:Z U175:C U175:B U175:A gnd gnds vdd vdds HS65_GSS_XNOR3X2
XU176 U176:Z U176:B U176:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU177 U177:Z U177:A gnd gnds vdd vdds HS65_GS_IVX9
XU178 U178:Z U178:A gnd gnds vdd vdds HS65_GS_IVX9
XU180 U180:Z U180:B U180:A gnd gnds vdd vdds HS65_GSS_XOR2X3
XU181 U181:Z U181:A gnd gnds vdd vdds HS65_GS_IVX9
XU182 U182:Z U182:A gnd gnds vdd vdds HS65_GS_IVX9
XU183 U183:Z U183:C U183:B U183:A gnd gnds vdd vdds HS65_GS_NOR3X4
XU184 U184:Z U184:C U184:B U184:A gnd gnds vdd vdds HS65_GS_NOR3AX2
XU185 U185:Z U185:A gnd gnds vdd vdds HS65_GS_IVX9
XU186 U186:Z U186:B U186:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU187 U187:Z U187:A gnd gnds vdd vdds HS65_GS_IVX9
XU188 U188:Z U188:B U188:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU189 U189:Z U189:B U189:A gnd gnds vdd vdds HS65_GS_NAND2AX7
XU190 U190:Z U190:C U190:B U190:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU191 U191:Z U191:B U191:A gnd gnds vdd vdds HS65_GSS_XNOR2X6
XU192 U192:Z U192:C U192:B U192:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU193 U193:Z U193:B U193:A gnd gnds vdd vdds HS65_GSS_XNOR2X6
XU194 U194:Z U194:C U194:B U194:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU195 U195:Z U195:B U195:A gnd gnds vdd vdds HS65_GSS_XNOR2X6
XU196 U196:Z U196:C U196:B U196:A gnd gnds vdd vdds HS65_GSS_XNOR3X2
XU197 U197:Z U197:B U197:A gnd gnds vdd vdds HS65_GSS_XNOR2X6
XU198 U198:Z U198:B U198:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU199 U199:Z U199:C U199:B U199:A gnd gnds vdd vdds HS65_GSS_XNOR3X2
XU200 U200:Z U200:B U200:A gnd gnds vdd vdds HS65_GSS_XNOR2X6
XU201 U201:Z U201:C U201:B U201:A gnd gnds vdd vdds HS65_GS_NAND3X5
XU202 U202:Z U202:C U202:B U202:A gnd gnds vdd vdds HS65_GS_NAND3X5
XU203 U203:Z U203:B U203:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU204 U204:Z U204:B U204:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU205 U205:Z U205:B U205:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU206 U206:Z U206:B U206:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU207 U207:Z U207:C U207:B U207:A gnd gnds vdd vdds HS65_GSS_XNOR3X2
XU208 U208:Z U208:B U208:A gnd gnds vdd vdds HS65_GSS_XNOR2X6
XU209 U209:Z U209:B U209:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU210 U210:Z U210:B U210:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU211 U211:Z U211:B U211:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU212 U212:Z U212:C U212:B U212:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU213 U213:Z U213:B U213:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU214 U214:Z U214:C U214:B U214:A gnd gnds vdd vdds HS65_GSS_XNOR3X2
XU215 U215:Z U215:B U215:A gnd gnds vdd vdds HS65_GSS_XNOR2X6
XU216 U216:Z U216:C U216:B U216:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU217 U217:Z U217:C U217:B U217:A gnd gnds vdd vdds HS65_GSS_XNOR3X2
XU218 U218:Z U218:B U218:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU219 U219:Z U219:B U219:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU220 U220:Z U220:C U220:B U220:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU221 U221:Z U221:C U221:B U221:A gnd gnds vdd vdds HS65_GSS_XNOR3X2
XU222 U222:Z U222:B U222:A gnd gnds vdd vdds HS65_GSS_XNOR2X6
XU223 U223:Z U223:B U223:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU224 U224:Z U224:B U224:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU225 U225:Z U225:B U225:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU226 U226:Z U226:B U226:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU227 U227:Z U227:B U227:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU228 U228:Z U228:B U228:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU229 U229:Z U229:B U229:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU230 U230:Z U230:B U230:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU231 U231:Z U231:B U231:A gnd gnds vdd vdds HS65_GS_NAND2X7
XU232 U232:Z U232:B U232:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU233 U233:Z U233:B U233:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU234 U234:Z U234:B U234:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU235 U235:Z U235:B U235:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU236 U236:Z U236:C U236:B U236:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU237 U237:Z U237:C U237:B U237:A gnd gnds vdd vdds HS65_GSS_XNOR3X2
XU238 U238:Z U238:B U238:A gnd gnds vdd vdds HS65_GSS_XNOR2X6
XU239 U239:Z U239:B U239:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU240 U240:Z U240:B U240:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU241 U241:Z U241:B U241:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU242 U242:Z U242:B U242:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU243 U243:Z U243:B U243:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU244 U244:Z U244:B U244:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU245 U245:Z U245:B U245:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU246 U246:Z U246:B U246:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU247 U247:Z U247:B U247:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU248 U248:Z U248:C U248:B U248:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU249 U249:Z U249:B U249:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU250 U250:Z U250:C U250:B U250:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU251 U251:Z U251:B U251:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU252 U252:Z U252:C U252:B U252:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU253 U253:Z U253:B U253:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU254 U254:Z U254:C U254:B U254:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU255 U255:Z U255:B U255:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU256 U256:Z U256:C U256:B U256:A gnd gnds vdd vdds HS65_GSS_XOR3X2
XU257 U257:Z U257:C U257:B U257:A gnd gnds vdd vdds HS65_GSS_XNOR3X2
XU258 U258:Z U258:B U258:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU259 U259:Z U259:B U259:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU260 U260:Z U260:B U260:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU261 U261:Z U261:B U261:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU262 U262:Z U262:B U262:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU263 U263:Z U263:B U263:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU264 U264:Z U264:B U264:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU265 U265:Z U265:B U265:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU266 U266:Z U266:B U266:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU267 U267:Z U267:B U267:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU268 U268:Z U268:B U268:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU269 U269:Z U269:B U269:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU270 U270:Z U270:B U270:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU271 U271:Z U271:B U271:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU272 U272:Z U272:B U272:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU273 U273:Z U273:B U273:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU274 U274:Z U274:B U274:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU275 U275:Z U275:B U275:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU276 U276:Z U276:B U276:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU277 U277:Z U277:B U277:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU278 U278:Z U278:B U278:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU279 U279:Z U279:B U279:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU280 U280:Z U280:B U280:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU281 U281:Z U281:B U281:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU282 U282:Z U282:B U282:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU283 U283:Z U283:B U283:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU284 U284:Z U284:B U284:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU285 U285:Z U285:B U285:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU286 U286:Z U286:B U286:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU287 U287:Z U287:B U287:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU288 U288:Z U288:B U288:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU289 U289:Z U289:B U289:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU290 U290:Z U290:B U290:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU291 U291:Z U291:B U291:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU292 U292:Z U292:B U292:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU293 U293:Z U293:B U293:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU294 U294:Z U294:B U294:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU295 U295:Z U295:B U295:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU296 U296:Z U296:B U296:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU297 U297:Z U297:B U297:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU298 U298:Z U298:B U298:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU299 U299:Z U299:B U299:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU300 U300:Z U300:B U300:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU301 U301:Z U301:B U301:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU302 U302:Z U302:B U302:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU303 U303:Z U303:B U303:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU304 U304:Z U304:B U304:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU305 U305:Z U305:B U305:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU306 U306:Z U306:B U306:A gnd gnds vdd vdds HS65_GSS_XOR2X6
XU307 U307:Z U307:B U307:A gnd gnds vdd vdds HS65_GS_NOR2X6
XU308 U308:Z U308:A gnd gnds vdd vdds HS65_GS_IVX9
XU309 U309:Z U309:A gnd gnds vdd vdds HS65_GS_IVX9
XU310 U310:Z U310:A gnd gnds vdd vdds HS65_GS_IVX9
XU311 U311:Z U311:A gnd gnds vdd vdds HS65_GS_IVX9
XU312 U312:Z U312:A gnd gnds vdd vdds HS65_GS_IVX9
XU313 U313:Z U313:A gnd gnds vdd vdds HS65_GS_IVX9
XU314 U314:Z U314:A gnd gnds vdd vdds HS65_GS_IVX9
XU315 U315:Z U315:B U315:A gnd gnds vdd vdds HS65_GSS_XNOR2X6
XU316 U316:Z U316:B U316:A gnd gnds vdd vdds HS65_GS_NOR2X6
.ENDS


******Simulation parameters*****

****Param definitions***
.param clk_period= '(1/500)*(0.000001)' 
+half_clk_period= '(clk_period/2)'
+double_clk_period= '(clk_period*2)'

.param fall_from_value=4e-09
+ fall_to_value=4.05e-09

.param init_delay = half_clk_period
+ rise_time= 50p
+ fall_time= 50p

**2.5 cycle simulation**
.param change_time='(half_clk_period/3)'
.param change_time_rise= '(change_time + 100ps)'
.param k_plus1= '(half_clk_period + change_time)'
.param k_plus1_rise = '(k_plus1 + 100ps)'
.param current_magnitude = 1.2mA
+rise_delay= 1.66344711153e-09s
+fall_delay= 'rise_delay+5p'
+rise_time_constant = 1ps
+fall_time_constant=130ps

.GLOBAL vdd gnd

Vvdd vdd 0 1
Vgnd agnd 0 0
Rgnd agnd gnd 0
VCk  clk   0  PULSE(0 1 init_delay rise_time fall_time half_clk_period clk_period)



******Instantiating the subckt*****

Xc499_clk_opFF
+ clk PNN1 PNN5 PNN9 PNN13 PNN17 PNN21 PNN25 PNN29 PNN33 
+ PNN37 PNN41 PNN45 PNN49 PNN53 PNN57 PNN61 PNN65 PNN69 PNN73 
+ PNN77 PNN81 PNN85 PNN89 PNN93 PNN97 PNN101 PNN105 PNN109 PNN113 
+ PNN117 PNN121 PNN125 PNN129 PNN130 PNN131 PNN132 PNN133 PNN134 PNN135 
+ PNN136 PNN137 Qout_PNN724 Qout_PNN725 Qout_PNN726 Qout_PNN727 Qout_PNN728 Qout_PNN729 Qout_PNN730 Qout_PNN731 
+ Qout_PNN732 Qout_PNN733 Qout_PNN734 Qout_PNN735 Qout_PNN736 Qout_PNN737 Qout_PNN738 Qout_PNN739 Qout_PNN740 Qout_PNN741 
+ Qout_PNN742 Qout_PNN743 Qout_PNN744 Qout_PNN745 Qout_PNN746 Qout_PNN747 Qout_PNN748 Qout_PNN749 Qout_PNN750 Qout_PNN751 
+ Qout_PNN752 Qout_PNN753 Qout_PNN754 Qout_PNN755  c499_clk_opFF

******Done instantiating the subckt*****


V1 PNN1 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V2 PNN5 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V3 PNN9 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V4 PNN13 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V5 PNN17 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V6 PNN21 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V7 PNN25 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V8 PNN29 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V9 PNN33 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V10 PNN37 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V11 PNN41 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V12 PNN45 0 PWL( 0  1 k_plus1 1 k_plus1_rise 0 5e-09 0)


V13 PNN49 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V14 PNN53 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V15 PNN57 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V16 PNN61 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V17 PNN65 0 PWL( 0  0 k_plus1 0 k_plus1_rise 1 5e-09 1)


V18 PNN69 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V19 PNN73 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V20 PNN77 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V21 PNN81 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V22 PNN85 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V23 PNN89 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V24 PNN93 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V25 PNN97 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V26 PNN101 0 PWL( 0  0 k_plus1 0 k_plus1_rise 1 5e-09 1)


V27 PNN105 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V28 PNN109 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V29 PNN113 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V30 PNN117 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V31 PNN121 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V32 PNN125 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V33 PNN129 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V34 PNN130 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V35 PNN131 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V36 PNN132 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V37 PNN133 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V38 PNN134 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V39 PNN135 0 PWL( 0  0 k_plus1 0 k_plus1_rise 0 5e-09 0)


V40 PNN136 0 PWL( 0  1 k_plus1 1 k_plus1_rise 1 5e-09 1)


V41 PNN137 0 PWL( 0  0 k_plus1 0 k_plus1_rise 1 5e-09 1)

**Initialising input of all FFs- commented this out. Doesnt help.PWL

**Initialising output of all FFs- trying..

**This is the initial value on the Qbar signal inside the DFF. 
.ic v(Xc499_clk_opFF.XiDFF_1_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_1_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_2_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_2_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_3_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_3_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_4_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_4_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_6_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_6_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_7_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_7_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_8_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_8_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_9_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_9_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_10_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_10_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_11_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_11_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_12_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_12_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_13_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_13_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_14_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_14_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_15_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_15_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_16_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_16_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_17_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_17_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_18_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_18_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_19_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_19_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_20_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_20_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_21_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_21_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_22_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_22_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_23_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_23_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_24_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_24_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_25_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_25_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_26_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_26_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_27_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_27_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_28_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_28_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_29_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_29_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_30_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_30_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_31_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_31_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_32_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_32_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_33_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_33_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_34_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_34_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_35_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_35_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_36_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_36_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_37_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_37_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_38_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_38_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_39_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_39_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_40_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XiDFF_40_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XiDFF_41_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XiDFF_41_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_1_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XoDFF_1_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XoDFF_2_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XoDFF_2_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XoDFF_3_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XoDFF_3_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XoDFF_4_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_4_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_5_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XoDFF_5_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XoDFF_6_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XoDFF_6_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XoDFF_7_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_7_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_8_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_8_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_9_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_9_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_10_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XoDFF_10_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XoDFF_11_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XoDFF_11_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XoDFF_12_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XoDFF_12_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XoDFF_13_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XoDFF_13_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XoDFF_14_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XoDFF_14_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XoDFF_15_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_15_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_16_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_16_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_17_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_17_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_18_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_18_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_19_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XoDFF_19_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XoDFF_20_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_20_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_21_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_21_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_22_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XoDFF_22_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XoDFF_23_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_23_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_24_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_24_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_25_q_reg.net0148:F59)= 0
.ic v(Xc499_clk_opFF.XoDFF_25_q_reg.net0148:F65)= 0

.ic v(Xc499_clk_opFF.XoDFF_26_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_26_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_27_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_27_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_28_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_28_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_29_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_29_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_30_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_30_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_31_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_31_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XoDFF_32_q_reg.net0148:F59)= 1
.ic v(Xc499_clk_opFF.XoDFF_32_q_reg.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG28_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG28_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG16_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG16_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG25_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG25_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG13_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG13_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG1_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG1_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG5_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG5_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG6_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG6_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG8_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG8_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG9_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG9_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG7_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG7_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG10_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG10_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG2_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG2_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG21_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG21_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG22_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG22_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG3_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG3_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG17_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG17_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG18_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG18_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG26_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG26_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG29_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG29_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG30_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG30_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG31_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG31_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG32_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG32_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG33_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG33_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG34_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG34_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG35_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG35_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG36_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG36_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG37_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG37_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG38_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG38_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG39_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG39_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG40_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG40_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG41_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG41_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG42_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG42_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG43_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG43_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG44_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG44_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG45_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG45_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG46_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG46_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG47_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG47_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG48_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG48_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG49_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG49_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG50_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG50_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG51_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG51_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG0_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG0_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG12_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG12_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG15_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG15_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG27_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG27_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG4_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG4_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG11_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG11_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG24_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG24_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG20_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG20_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG23_S2.net0148:F59)= 0
.ic v(Xc499_clk_opFF.Xclk_r_REG23_S2.net0148:F65)= 0

.ic v(Xc499_clk_opFF.Xclk_r_REG19_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG19_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.Xclk_r_REG14_S2.net0148:F59)= 1
.ic v(Xc499_clk_opFF.Xclk_r_REG14_S2.net0148:F65)= 1

.ic v(Xc499_clk_opFF.XiDFF_5_q_reg.net0139:F125)= 1



**Initialising primary outputs to 0..commented out right now



.control
option rshunt = 1e12
option itl4 = 100  reltol =0.005  trtol=8 pivtol=1e-11  abstol=1e-10 
**option CONVERGE=-1
tran 20ps 5e-09s

**Uncomment the following and run this spice file, if you need a waveform
**write waveform_file.raw v(clk) v(input_dec_2_) v(input_dec_1_) v(input_dec_0_)  v(output_dec_3_) v(output_dec_1_) 
*+v.xdecoder_behav_pnr.xu11.vcharge#branch 



**************************** Measuring Flip Flop output at 2nd falling edge *************************************************
meas tran ff_op_fall_0 MAX v(Xc499_clk_opFF.iDFF_1_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_1 MAX v(Xc499_clk_opFF.iDFF_2_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_2 MAX v(Xc499_clk_opFF.iDFF_3_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_3 MAX v(Xc499_clk_opFF.iDFF_4_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_4 MAX v(Xc499_clk_opFF.iDFF_6_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_5 MAX v(Xc499_clk_opFF.iDFF_7_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_6 MAX v(Xc499_clk_opFF.iDFF_8_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_7 MAX v(Xc499_clk_opFF.iDFF_9_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_8 MAX v(Xc499_clk_opFF.iDFF_10_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_9 MAX v(Xc499_clk_opFF.iDFF_11_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_10 MAX v(Xc499_clk_opFF.iDFF_12_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_11 MAX v(Xc499_clk_opFF.iDFF_13_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_12 MAX v(Xc499_clk_opFF.iDFF_14_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_13 MAX v(Xc499_clk_opFF.iDFF_15_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_14 MAX v(Xc499_clk_opFF.iDFF_16_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_15 MAX v(Xc499_clk_opFF.iDFF_17_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_16 MAX v(Xc499_clk_opFF.iDFF_18_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_17 MAX v(Xc499_clk_opFF.iDFF_19_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_18 MAX v(Xc499_clk_opFF.iDFF_20_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_19 MAX v(Xc499_clk_opFF.iDFF_21_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_20 MAX v(Xc499_clk_opFF.iDFF_22_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_21 MAX v(Xc499_clk_opFF.iDFF_23_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_22 MAX v(Xc499_clk_opFF.iDFF_24_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_23 MAX v(Xc499_clk_opFF.iDFF_25_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_24 MAX v(Xc499_clk_opFF.iDFF_26_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_25 MAX v(Xc499_clk_opFF.iDFF_27_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_26 MAX v(Xc499_clk_opFF.iDFF_28_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_27 MAX v(Xc499_clk_opFF.iDFF_29_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_28 MAX v(Xc499_clk_opFF.iDFF_30_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_29 MAX v(Xc499_clk_opFF.iDFF_31_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_30 MAX v(Xc499_clk_opFF.iDFF_32_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_31 MAX v(Xc499_clk_opFF.iDFF_33_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_32 MAX v(Xc499_clk_opFF.iDFF_34_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_33 MAX v(Xc499_clk_opFF.iDFF_35_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_34 MAX v(Xc499_clk_opFF.iDFF_36_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_35 MAX v(Xc499_clk_opFF.iDFF_37_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_36 MAX v(Xc499_clk_opFF.iDFF_38_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_37 MAX v(Xc499_clk_opFF.iDFF_39_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_38 MAX v(Xc499_clk_opFF.iDFF_40_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_39 MAX v(Xc499_clk_opFF.iDFF_41_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_40 MAX v(Xc499_clk_opFF.oDFF_1_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_41 MAX v(Xc499_clk_opFF.oDFF_2_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_42 MAX v(Xc499_clk_opFF.oDFF_3_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_43 MAX v(Xc499_clk_opFF.oDFF_4_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_44 MAX v(Xc499_clk_opFF.oDFF_5_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_45 MAX v(Xc499_clk_opFF.oDFF_6_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_46 MAX v(Xc499_clk_opFF.oDFF_7_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_47 MAX v(Xc499_clk_opFF.oDFF_8_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_48 MAX v(Xc499_clk_opFF.oDFF_9_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_49 MAX v(Xc499_clk_opFF.oDFF_10_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_50 MAX v(Xc499_clk_opFF.oDFF_11_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_51 MAX v(Xc499_clk_opFF.oDFF_12_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_52 MAX v(Xc499_clk_opFF.oDFF_13_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_53 MAX v(Xc499_clk_opFF.oDFF_14_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_54 MAX v(Xc499_clk_opFF.oDFF_15_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_55 MAX v(Xc499_clk_opFF.oDFF_16_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_56 MAX v(Xc499_clk_opFF.oDFF_17_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_57 MAX v(Xc499_clk_opFF.oDFF_18_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_58 MAX v(Xc499_clk_opFF.oDFF_19_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_59 MAX v(Xc499_clk_opFF.oDFF_20_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_60 MAX v(Xc499_clk_opFF.oDFF_21_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_61 MAX v(Xc499_clk_opFF.oDFF_22_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_62 MAX v(Xc499_clk_opFF.oDFF_23_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_63 MAX v(Xc499_clk_opFF.oDFF_24_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_64 MAX v(Xc499_clk_opFF.oDFF_25_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_65 MAX v(Xc499_clk_opFF.oDFF_26_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_66 MAX v(Xc499_clk_opFF.oDFF_27_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_67 MAX v(Xc499_clk_opFF.oDFF_28_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_68 MAX v(Xc499_clk_opFF.oDFF_29_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_69 MAX v(Xc499_clk_opFF.oDFF_30_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_70 MAX v(Xc499_clk_opFF.oDFF_31_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_71 MAX v(Xc499_clk_opFF.oDFF_32_q_reg:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_72 MAX v(Xc499_clk_opFF.clk_r_REG28_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_73 MAX v(Xc499_clk_opFF.clk_r_REG16_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_74 MAX v(Xc499_clk_opFF.clk_r_REG25_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_75 MAX v(Xc499_clk_opFF.clk_r_REG13_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_76 MAX v(Xc499_clk_opFF.clk_r_REG1_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_77 MAX v(Xc499_clk_opFF.clk_r_REG5_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_78 MAX v(Xc499_clk_opFF.clk_r_REG6_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_79 MAX v(Xc499_clk_opFF.clk_r_REG8_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_80 MAX v(Xc499_clk_opFF.clk_r_REG9_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_81 MAX v(Xc499_clk_opFF.clk_r_REG7_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_82 MAX v(Xc499_clk_opFF.clk_r_REG10_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_83 MAX v(Xc499_clk_opFF.clk_r_REG2_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_84 MAX v(Xc499_clk_opFF.clk_r_REG21_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_85 MAX v(Xc499_clk_opFF.clk_r_REG22_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_86 MAX v(Xc499_clk_opFF.clk_r_REG3_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_87 MAX v(Xc499_clk_opFF.clk_r_REG17_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_88 MAX v(Xc499_clk_opFF.clk_r_REG18_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_89 MAX v(Xc499_clk_opFF.clk_r_REG26_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_90 MAX v(Xc499_clk_opFF.clk_r_REG29_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_91 MAX v(Xc499_clk_opFF.clk_r_REG30_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_92 MAX v(Xc499_clk_opFF.clk_r_REG31_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_93 MAX v(Xc499_clk_opFF.clk_r_REG32_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_94 MAX v(Xc499_clk_opFF.clk_r_REG33_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_95 MAX v(Xc499_clk_opFF.clk_r_REG34_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_96 MAX v(Xc499_clk_opFF.clk_r_REG35_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_97 MAX v(Xc499_clk_opFF.clk_r_REG36_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_98 MAX v(Xc499_clk_opFF.clk_r_REG37_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_99 MAX v(Xc499_clk_opFF.clk_r_REG38_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_100 MAX v(Xc499_clk_opFF.clk_r_REG39_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_101 MAX v(Xc499_clk_opFF.clk_r_REG40_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_102 MAX v(Xc499_clk_opFF.clk_r_REG41_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_103 MAX v(Xc499_clk_opFF.clk_r_REG42_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_104 MAX v(Xc499_clk_opFF.clk_r_REG43_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_105 MAX v(Xc499_clk_opFF.clk_r_REG44_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_106 MAX v(Xc499_clk_opFF.clk_r_REG45_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_107 MAX v(Xc499_clk_opFF.clk_r_REG46_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_108 MAX v(Xc499_clk_opFF.clk_r_REG47_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_109 MAX v(Xc499_clk_opFF.clk_r_REG48_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_110 MAX v(Xc499_clk_opFF.clk_r_REG49_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_111 MAX v(Xc499_clk_opFF.clk_r_REG50_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_112 MAX v(Xc499_clk_opFF.clk_r_REG51_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_113 MAX v(Xc499_clk_opFF.clk_r_REG0_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_114 MAX v(Xc499_clk_opFF.clk_r_REG12_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_115 MAX v(Xc499_clk_opFF.clk_r_REG15_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_116 MAX v(Xc499_clk_opFF.clk_r_REG27_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_117 MAX v(Xc499_clk_opFF.clk_r_REG4_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_118 MAX v(Xc499_clk_opFF.clk_r_REG11_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_119 MAX v(Xc499_clk_opFF.clk_r_REG24_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_120 MAX v(Xc499_clk_opFF.clk_r_REG20_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_121 MAX v(Xc499_clk_opFF.clk_r_REG23_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_122 MAX v(Xc499_clk_opFF.clk_r_REG19_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_123 MAX v(Xc499_clk_opFF.clk_r_REG14_S2:Q) from=4e-09s to=4.05e-09s
meas tran ff_op_fall_124 MAX v(Xc499_clk_opFF.iDFF_5_q_reg:QN) from=4e-09s to=4.05e-09s


**************************** Measuring Flip Flop output at 2nd rising edge *************************************************
meas tran ff_op_rise_0 MAX v(Xc499_clk_opFF.iDFF_1_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_1 MAX v(Xc499_clk_opFF.iDFF_2_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_2 MAX v(Xc499_clk_opFF.iDFF_3_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_3 MAX v(Xc499_clk_opFF.iDFF_4_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_4 MAX v(Xc499_clk_opFF.iDFF_6_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_5 MAX v(Xc499_clk_opFF.iDFF_7_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_6 MAX v(Xc499_clk_opFF.iDFF_8_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_7 MAX v(Xc499_clk_opFF.iDFF_9_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_8 MAX v(Xc499_clk_opFF.iDFF_10_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_9 MAX v(Xc499_clk_opFF.iDFF_11_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_10 MAX v(Xc499_clk_opFF.iDFF_12_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_11 MAX v(Xc499_clk_opFF.iDFF_13_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_12 MAX v(Xc499_clk_opFF.iDFF_14_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_13 MAX v(Xc499_clk_opFF.iDFF_15_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_14 MAX v(Xc499_clk_opFF.iDFF_16_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_15 MAX v(Xc499_clk_opFF.iDFF_17_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_16 MAX v(Xc499_clk_opFF.iDFF_18_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_17 MAX v(Xc499_clk_opFF.iDFF_19_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_18 MAX v(Xc499_clk_opFF.iDFF_20_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_19 MAX v(Xc499_clk_opFF.iDFF_21_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_20 MAX v(Xc499_clk_opFF.iDFF_22_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_21 MAX v(Xc499_clk_opFF.iDFF_23_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_22 MAX v(Xc499_clk_opFF.iDFF_24_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_23 MAX v(Xc499_clk_opFF.iDFF_25_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_24 MAX v(Xc499_clk_opFF.iDFF_26_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_25 MAX v(Xc499_clk_opFF.iDFF_27_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_26 MAX v(Xc499_clk_opFF.iDFF_28_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_27 MAX v(Xc499_clk_opFF.iDFF_29_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_28 MAX v(Xc499_clk_opFF.iDFF_30_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_29 MAX v(Xc499_clk_opFF.iDFF_31_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_30 MAX v(Xc499_clk_opFF.iDFF_32_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_31 MAX v(Xc499_clk_opFF.iDFF_33_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_32 MAX v(Xc499_clk_opFF.iDFF_34_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_33 MAX v(Xc499_clk_opFF.iDFF_35_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_34 MAX v(Xc499_clk_opFF.iDFF_36_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_35 MAX v(Xc499_clk_opFF.iDFF_37_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_36 MAX v(Xc499_clk_opFF.iDFF_38_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_37 MAX v(Xc499_clk_opFF.iDFF_39_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_38 MAX v(Xc499_clk_opFF.iDFF_40_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_39 MAX v(Xc499_clk_opFF.iDFF_41_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_40 MAX v(Xc499_clk_opFF.oDFF_1_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_41 MAX v(Xc499_clk_opFF.oDFF_2_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_42 MAX v(Xc499_clk_opFF.oDFF_3_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_43 MAX v(Xc499_clk_opFF.oDFF_4_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_44 MAX v(Xc499_clk_opFF.oDFF_5_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_45 MAX v(Xc499_clk_opFF.oDFF_6_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_46 MAX v(Xc499_clk_opFF.oDFF_7_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_47 MAX v(Xc499_clk_opFF.oDFF_8_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_48 MAX v(Xc499_clk_opFF.oDFF_9_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_49 MAX v(Xc499_clk_opFF.oDFF_10_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_50 MAX v(Xc499_clk_opFF.oDFF_11_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_51 MAX v(Xc499_clk_opFF.oDFF_12_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_52 MAX v(Xc499_clk_opFF.oDFF_13_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_53 MAX v(Xc499_clk_opFF.oDFF_14_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_54 MAX v(Xc499_clk_opFF.oDFF_15_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_55 MAX v(Xc499_clk_opFF.oDFF_16_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_56 MAX v(Xc499_clk_opFF.oDFF_17_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_57 MAX v(Xc499_clk_opFF.oDFF_18_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_58 MAX v(Xc499_clk_opFF.oDFF_19_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_59 MAX v(Xc499_clk_opFF.oDFF_20_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_60 MAX v(Xc499_clk_opFF.oDFF_21_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_61 MAX v(Xc499_clk_opFF.oDFF_22_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_62 MAX v(Xc499_clk_opFF.oDFF_23_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_63 MAX v(Xc499_clk_opFF.oDFF_24_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_64 MAX v(Xc499_clk_opFF.oDFF_25_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_65 MAX v(Xc499_clk_opFF.oDFF_26_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_66 MAX v(Xc499_clk_opFF.oDFF_27_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_67 MAX v(Xc499_clk_opFF.oDFF_28_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_68 MAX v(Xc499_clk_opFF.oDFF_29_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_69 MAX v(Xc499_clk_opFF.oDFF_30_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_70 MAX v(Xc499_clk_opFF.oDFF_31_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_71 MAX v(Xc499_clk_opFF.oDFF_32_q_reg:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_72 MAX v(Xc499_clk_opFF.clk_r_REG28_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_73 MAX v(Xc499_clk_opFF.clk_r_REG16_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_74 MAX v(Xc499_clk_opFF.clk_r_REG25_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_75 MAX v(Xc499_clk_opFF.clk_r_REG13_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_76 MAX v(Xc499_clk_opFF.clk_r_REG1_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_77 MAX v(Xc499_clk_opFF.clk_r_REG5_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_78 MAX v(Xc499_clk_opFF.clk_r_REG6_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_79 MAX v(Xc499_clk_opFF.clk_r_REG8_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_80 MAX v(Xc499_clk_opFF.clk_r_REG9_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_81 MAX v(Xc499_clk_opFF.clk_r_REG7_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_82 MAX v(Xc499_clk_opFF.clk_r_REG10_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_83 MAX v(Xc499_clk_opFF.clk_r_REG2_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_84 MAX v(Xc499_clk_opFF.clk_r_REG21_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_85 MAX v(Xc499_clk_opFF.clk_r_REG22_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_86 MAX v(Xc499_clk_opFF.clk_r_REG3_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_87 MAX v(Xc499_clk_opFF.clk_r_REG17_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_88 MAX v(Xc499_clk_opFF.clk_r_REG18_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_89 MAX v(Xc499_clk_opFF.clk_r_REG26_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_90 MAX v(Xc499_clk_opFF.clk_r_REG29_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_91 MAX v(Xc499_clk_opFF.clk_r_REG30_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_92 MAX v(Xc499_clk_opFF.clk_r_REG31_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_93 MAX v(Xc499_clk_opFF.clk_r_REG32_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_94 MAX v(Xc499_clk_opFF.clk_r_REG33_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_95 MAX v(Xc499_clk_opFF.clk_r_REG34_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_96 MAX v(Xc499_clk_opFF.clk_r_REG35_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_97 MAX v(Xc499_clk_opFF.clk_r_REG36_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_98 MAX v(Xc499_clk_opFF.clk_r_REG37_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_99 MAX v(Xc499_clk_opFF.clk_r_REG38_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_100 MAX v(Xc499_clk_opFF.clk_r_REG39_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_101 MAX v(Xc499_clk_opFF.clk_r_REG40_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_102 MAX v(Xc499_clk_opFF.clk_r_REG41_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_103 MAX v(Xc499_clk_opFF.clk_r_REG42_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_104 MAX v(Xc499_clk_opFF.clk_r_REG43_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_105 MAX v(Xc499_clk_opFF.clk_r_REG44_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_106 MAX v(Xc499_clk_opFF.clk_r_REG45_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_107 MAX v(Xc499_clk_opFF.clk_r_REG46_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_108 MAX v(Xc499_clk_opFF.clk_r_REG47_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_109 MAX v(Xc499_clk_opFF.clk_r_REG48_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_110 MAX v(Xc499_clk_opFF.clk_r_REG49_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_111 MAX v(Xc499_clk_opFF.clk_r_REG50_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_112 MAX v(Xc499_clk_opFF.clk_r_REG51_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_113 MAX v(Xc499_clk_opFF.clk_r_REG0_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_114 MAX v(Xc499_clk_opFF.clk_r_REG12_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_115 MAX v(Xc499_clk_opFF.clk_r_REG15_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_116 MAX v(Xc499_clk_opFF.clk_r_REG27_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_117 MAX v(Xc499_clk_opFF.clk_r_REG4_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_118 MAX v(Xc499_clk_opFF.clk_r_REG11_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_119 MAX v(Xc499_clk_opFF.clk_r_REG24_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_120 MAX v(Xc499_clk_opFF.clk_r_REG20_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_121 MAX v(Xc499_clk_opFF.clk_r_REG23_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_122 MAX v(Xc499_clk_opFF.clk_r_REG19_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_123 MAX v(Xc499_clk_opFF.clk_r_REG14_S2:Q) from=3e-09s to=3.05e-09s
meas tran ff_op_rise_124 MAX v(Xc499_clk_opFF.iDFF_5_q_reg:QN) from=3e-09s to=3.05e-09s


**************************** Measuring Flip Flop output t=0 *************************************************
meas tran ff_op_time0_0 MAX v(Xc499_clk_opFF.iDFF_1_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_1 MAX v(Xc499_clk_opFF.iDFF_2_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_2 MAX v(Xc499_clk_opFF.iDFF_3_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_3 MAX v(Xc499_clk_opFF.iDFF_4_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_4 MAX v(Xc499_clk_opFF.iDFF_6_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_5 MAX v(Xc499_clk_opFF.iDFF_7_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_6 MAX v(Xc499_clk_opFF.iDFF_8_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_7 MAX v(Xc499_clk_opFF.iDFF_9_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_8 MAX v(Xc499_clk_opFF.iDFF_10_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_9 MAX v(Xc499_clk_opFF.iDFF_11_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_10 MAX v(Xc499_clk_opFF.iDFF_12_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_11 MAX v(Xc499_clk_opFF.iDFF_13_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_12 MAX v(Xc499_clk_opFF.iDFF_14_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_13 MAX v(Xc499_clk_opFF.iDFF_15_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_14 MAX v(Xc499_clk_opFF.iDFF_16_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_15 MAX v(Xc499_clk_opFF.iDFF_17_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_16 MAX v(Xc499_clk_opFF.iDFF_18_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_17 MAX v(Xc499_clk_opFF.iDFF_19_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_18 MAX v(Xc499_clk_opFF.iDFF_20_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_19 MAX v(Xc499_clk_opFF.iDFF_21_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_20 MAX v(Xc499_clk_opFF.iDFF_22_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_21 MAX v(Xc499_clk_opFF.iDFF_23_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_22 MAX v(Xc499_clk_opFF.iDFF_24_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_23 MAX v(Xc499_clk_opFF.iDFF_25_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_24 MAX v(Xc499_clk_opFF.iDFF_26_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_25 MAX v(Xc499_clk_opFF.iDFF_27_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_26 MAX v(Xc499_clk_opFF.iDFF_28_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_27 MAX v(Xc499_clk_opFF.iDFF_29_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_28 MAX v(Xc499_clk_opFF.iDFF_30_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_29 MAX v(Xc499_clk_opFF.iDFF_31_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_30 MAX v(Xc499_clk_opFF.iDFF_32_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_31 MAX v(Xc499_clk_opFF.iDFF_33_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_32 MAX v(Xc499_clk_opFF.iDFF_34_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_33 MAX v(Xc499_clk_opFF.iDFF_35_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_34 MAX v(Xc499_clk_opFF.iDFF_36_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_35 MAX v(Xc499_clk_opFF.iDFF_37_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_36 MAX v(Xc499_clk_opFF.iDFF_38_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_37 MAX v(Xc499_clk_opFF.iDFF_39_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_38 MAX v(Xc499_clk_opFF.iDFF_40_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_39 MAX v(Xc499_clk_opFF.iDFF_41_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_40 MAX v(Xc499_clk_opFF.oDFF_1_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_41 MAX v(Xc499_clk_opFF.oDFF_2_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_42 MAX v(Xc499_clk_opFF.oDFF_3_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_43 MAX v(Xc499_clk_opFF.oDFF_4_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_44 MAX v(Xc499_clk_opFF.oDFF_5_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_45 MAX v(Xc499_clk_opFF.oDFF_6_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_46 MAX v(Xc499_clk_opFF.oDFF_7_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_47 MAX v(Xc499_clk_opFF.oDFF_8_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_48 MAX v(Xc499_clk_opFF.oDFF_9_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_49 MAX v(Xc499_clk_opFF.oDFF_10_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_50 MAX v(Xc499_clk_opFF.oDFF_11_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_51 MAX v(Xc499_clk_opFF.oDFF_12_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_52 MAX v(Xc499_clk_opFF.oDFF_13_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_53 MAX v(Xc499_clk_opFF.oDFF_14_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_54 MAX v(Xc499_clk_opFF.oDFF_15_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_55 MAX v(Xc499_clk_opFF.oDFF_16_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_56 MAX v(Xc499_clk_opFF.oDFF_17_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_57 MAX v(Xc499_clk_opFF.oDFF_18_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_58 MAX v(Xc499_clk_opFF.oDFF_19_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_59 MAX v(Xc499_clk_opFF.oDFF_20_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_60 MAX v(Xc499_clk_opFF.oDFF_21_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_61 MAX v(Xc499_clk_opFF.oDFF_22_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_62 MAX v(Xc499_clk_opFF.oDFF_23_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_63 MAX v(Xc499_clk_opFF.oDFF_24_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_64 MAX v(Xc499_clk_opFF.oDFF_25_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_65 MAX v(Xc499_clk_opFF.oDFF_26_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_66 MAX v(Xc499_clk_opFF.oDFF_27_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_67 MAX v(Xc499_clk_opFF.oDFF_28_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_68 MAX v(Xc499_clk_opFF.oDFF_29_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_69 MAX v(Xc499_clk_opFF.oDFF_30_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_70 MAX v(Xc499_clk_opFF.oDFF_31_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_71 MAX v(Xc499_clk_opFF.oDFF_32_q_reg:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_72 MAX v(Xc499_clk_opFF.clk_r_REG28_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_73 MAX v(Xc499_clk_opFF.clk_r_REG16_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_74 MAX v(Xc499_clk_opFF.clk_r_REG25_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_75 MAX v(Xc499_clk_opFF.clk_r_REG13_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_76 MAX v(Xc499_clk_opFF.clk_r_REG1_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_77 MAX v(Xc499_clk_opFF.clk_r_REG5_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_78 MAX v(Xc499_clk_opFF.clk_r_REG6_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_79 MAX v(Xc499_clk_opFF.clk_r_REG8_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_80 MAX v(Xc499_clk_opFF.clk_r_REG9_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_81 MAX v(Xc499_clk_opFF.clk_r_REG7_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_82 MAX v(Xc499_clk_opFF.clk_r_REG10_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_83 MAX v(Xc499_clk_opFF.clk_r_REG2_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_84 MAX v(Xc499_clk_opFF.clk_r_REG21_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_85 MAX v(Xc499_clk_opFF.clk_r_REG22_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_86 MAX v(Xc499_clk_opFF.clk_r_REG3_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_87 MAX v(Xc499_clk_opFF.clk_r_REG17_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_88 MAX v(Xc499_clk_opFF.clk_r_REG18_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_89 MAX v(Xc499_clk_opFF.clk_r_REG26_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_90 MAX v(Xc499_clk_opFF.clk_r_REG29_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_91 MAX v(Xc499_clk_opFF.clk_r_REG30_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_92 MAX v(Xc499_clk_opFF.clk_r_REG31_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_93 MAX v(Xc499_clk_opFF.clk_r_REG32_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_94 MAX v(Xc499_clk_opFF.clk_r_REG33_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_95 MAX v(Xc499_clk_opFF.clk_r_REG34_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_96 MAX v(Xc499_clk_opFF.clk_r_REG35_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_97 MAX v(Xc499_clk_opFF.clk_r_REG36_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_98 MAX v(Xc499_clk_opFF.clk_r_REG37_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_99 MAX v(Xc499_clk_opFF.clk_r_REG38_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_100 MAX v(Xc499_clk_opFF.clk_r_REG39_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_101 MAX v(Xc499_clk_opFF.clk_r_REG40_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_102 MAX v(Xc499_clk_opFF.clk_r_REG41_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_103 MAX v(Xc499_clk_opFF.clk_r_REG42_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_104 MAX v(Xc499_clk_opFF.clk_r_REG43_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_105 MAX v(Xc499_clk_opFF.clk_r_REG44_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_106 MAX v(Xc499_clk_opFF.clk_r_REG45_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_107 MAX v(Xc499_clk_opFF.clk_r_REG46_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_108 MAX v(Xc499_clk_opFF.clk_r_REG47_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_109 MAX v(Xc499_clk_opFF.clk_r_REG48_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_110 MAX v(Xc499_clk_opFF.clk_r_REG49_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_111 MAX v(Xc499_clk_opFF.clk_r_REG50_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_112 MAX v(Xc499_clk_opFF.clk_r_REG51_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_113 MAX v(Xc499_clk_opFF.clk_r_REG0_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_114 MAX v(Xc499_clk_opFF.clk_r_REG12_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_115 MAX v(Xc499_clk_opFF.clk_r_REG15_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_116 MAX v(Xc499_clk_opFF.clk_r_REG27_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_117 MAX v(Xc499_clk_opFF.clk_r_REG4_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_118 MAX v(Xc499_clk_opFF.clk_r_REG11_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_119 MAX v(Xc499_clk_opFF.clk_r_REG24_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_120 MAX v(Xc499_clk_opFF.clk_r_REG20_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_121 MAX v(Xc499_clk_opFF.clk_r_REG23_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_122 MAX v(Xc499_clk_opFF.clk_r_REG19_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_123 MAX v(Xc499_clk_opFF.clk_r_REG14_S2:Q) from=0.01e-9s to=0.05e-9s
meas tran ff_op_time0_124 MAX v(Xc499_clk_opFF.iDFF_5_q_reg:QN) from=0.01e-9s to=0.05e-9s


***************** saving the outputs at the 2nd falling edge ****************
echo "$&ff_op_fall_0" , > glitch_report_outputs_1.csv  $$New file
echo "$&ff_op_fall_1" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_2" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_3" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_4" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_5" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_6" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_7" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_8" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_9" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_10" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_11" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_12" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_13" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_14" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_15" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_16" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_17" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_18" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_19" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_20" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_21" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_22" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_23" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_24" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_25" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_26" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_27" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_28" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_29" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_30" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_31" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_32" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_33" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_34" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_35" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_36" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_37" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_38" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_39" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_40" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_41" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_42" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_43" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_44" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_45" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_46" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_47" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_48" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_49" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_50" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_51" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_52" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_53" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_54" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_55" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_56" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_57" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_58" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_59" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_60" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_61" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_62" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_63" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_64" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_65" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_66" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_67" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_68" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_69" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_70" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_71" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_72" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_73" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_74" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_75" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_76" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_77" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_78" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_79" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_80" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_81" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_82" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_83" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_84" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_85" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_86" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_87" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_88" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_89" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_90" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_91" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_92" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_93" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_94" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_95" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_96" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_97" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_98" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_99" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_100" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_101" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_102" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_103" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_104" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_105" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_106" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_107" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_108" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_109" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_110" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_111" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_112" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_113" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_114" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_115" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_116" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_117" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_118" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_119" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_120" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_121" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_122" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_123" , >> glitch_report_outputs_1.csv  $$Appending to the file
echo "$&ff_op_fall_124" , >> glitch_report_outputs_1.csv  $$Appending to the file


***************** saving the outputs at the 2nd rising edge ****************
echo "$&ff_op_rise_0" , > glitch_report_outputs_rise_1.csv  $$New file
echo "$&ff_op_rise_1" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_2" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_3" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_4" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_5" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_6" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_7" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_8" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_9" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_10" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_11" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_12" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_13" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_14" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_15" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_16" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_17" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_18" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_19" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_20" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_21" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_22" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_23" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_24" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_25" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_26" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_27" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_28" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_29" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_30" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_31" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_32" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_33" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_34" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_35" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_36" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_37" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_38" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_39" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_40" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_41" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_42" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_43" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_44" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_45" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_46" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_47" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_48" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_49" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_50" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_51" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_52" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_53" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_54" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_55" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_56" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_57" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_58" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_59" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_60" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_61" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_62" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_63" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_64" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_65" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_66" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_67" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_68" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_69" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_70" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_71" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_72" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_73" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_74" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_75" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_76" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_77" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_78" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_79" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_80" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_81" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_82" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_83" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_84" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_85" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_86" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_87" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_88" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_89" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_90" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_91" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_92" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_93" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_94" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_95" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_96" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_97" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_98" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_99" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_100" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_101" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_102" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_103" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_104" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_105" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_106" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_107" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_108" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_109" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_110" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_111" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_112" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_113" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_114" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_115" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_116" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_117" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_118" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_119" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_120" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_121" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_122" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_123" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file
echo "$&ff_op_rise_124" , >> glitch_report_outputs_rise_1.csv  $$Appending to the file


***************** saving the outputs at time=0 ****************
echo "$&ff_op_time0_0" , > glitch_report_outputs_time0_1.csv  $$New file
echo "$&ff_op_time0_1" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_2" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_3" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_4" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_5" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_6" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_7" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_8" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_9" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_10" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_11" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_12" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_13" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_14" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_15" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_16" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_17" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_18" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_19" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_20" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_21" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_22" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_23" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_24" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_25" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_26" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_27" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_28" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_29" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_30" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_31" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_32" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_33" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_34" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_35" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_36" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_37" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_38" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_39" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_40" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_41" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_42" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_43" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_44" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_45" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_46" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_47" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_48" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_49" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_50" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_51" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_52" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_53" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_54" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_55" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_56" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_57" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_58" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_59" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_60" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_61" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_62" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_63" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_64" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_65" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_66" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_67" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_68" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_69" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_70" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_71" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_72" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_73" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_74" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_75" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_76" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_77" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_78" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_79" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_80" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_81" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_82" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_83" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_84" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_85" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_86" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_87" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_88" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_89" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_90" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_91" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_92" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_93" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_94" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_95" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_96" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_97" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_98" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_99" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_100" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_101" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_102" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_103" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_104" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_105" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_106" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_107" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_108" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_109" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_110" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_111" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_112" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_113" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_114" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_115" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_116" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_117" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_118" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_119" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_120" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_121" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_122" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_123" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file
echo "$&ff_op_time0_124" , >> glitch_report_outputs_time0_1.csv  $$Appending to the file

quit

.endc


.end

** NUMBER OF OUTPUT PINS = 125
