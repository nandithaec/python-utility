********** Glitched induced version of LIBRARY : test_lib.sp **********



******************************* ORIGINAL SUBCIRCUIT : HS65_GS_AO212X4 ******************************* 

.SUBCKT HS65_GS_AO212X4 Z E D C B A gnd gnd vdd vdd
*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4

****** HS65_GS_AO212X4 : Glitched version 1 : glitch at net044:F64 ******

.SUBCKT HS65_GS_AO212X4_1 Z E D C B A gnd gnd vdd vdd
**PMOS current injection
Icharge 0 net044:F64 EXP (0 current_magnitude/3 rise_delay rise_time_constant fall_delay fall_time_constant)

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4_1

****** HS65_GS_AO212X4 : Glitched version 2 : glitch at net029:F50 ******

.SUBCKT HS65_GS_AO212X4_2 Z E D C B A gnd gnd vdd vdd
**PMOS current injection
Icharge 0 net029:F50 EXP (0 current_magnitude/3 rise_delay rise_time_constant fall_delay fall_time_constant)

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4_2

****** HS65_GS_AO212X4 : Glitched version 3 : glitch at net029:F42 ******

.SUBCKT HS65_GS_AO212X4_3 Z E D C B A gnd gnd vdd vdd
**NMOS current injection
Icharge net029:F42 0 EXP (0 current_magnitude rise_delay rise_time_constant fall_delay fall_time_constant)

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4_3

****** HS65_GS_AO212X4 : Glitched version 4 : glitch at net029:F36 ******

.SUBCKT HS65_GS_AO212X4_4 Z E D C B A gnd gnd vdd vdd
**NMOS current injection
Icharge net029:F36 0 EXP (0 current_magnitude rise_delay rise_time_constant fall_delay fall_time_constant)

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4_4

****** HS65_GS_AO212X4 : Glitched version 5 : glitch at net029:F60 ******

.SUBCKT HS65_GS_AO212X4_5 Z E D C B A gnd gnd vdd vdd
**PMOS current injection
Icharge 0 net029:F60 EXP (0 current_magnitude/3 rise_delay rise_time_constant fall_delay fall_time_constant)

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4_5

****** HS65_GS_AO212X4 : Glitched version 6 : glitch at Z:F24 ******

.SUBCKT HS65_GS_AO212X4_6 Z E D C B A gnd gnd vdd vdd
**NMOS current injection
Icharge Z:F24 0 EXP (0 current_magnitude rise_delay rise_time_constant fall_delay fall_time_constant)

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4_6

****** HS65_GS_AO212X4 : Glitched version 7 : glitch at net040:F70 ******

.SUBCKT HS65_GS_AO212X4_7 Z E D C B A gnd gnd vdd vdd
**PMOS current injection
Icharge 0 net040:F70 EXP (0 current_magnitude/3 rise_delay rise_time_constant fall_delay fall_time_constant)

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4_7

****** HS65_GS_AO212X4 : Glitched version 8 : glitch at net040:F68 ******

.SUBCKT HS65_GS_AO212X4_8 Z E D C B A gnd gnd vdd vdd
**PMOS current injection
Icharge 0 net040:F68 EXP (0 current_magnitude/3 rise_delay rise_time_constant fall_delay fall_time_constant)

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4_8

****** HS65_GS_AO212X4 : Glitched version 9 : glitch at Z:F46 ******

.SUBCKT HS65_GS_AO212X4_9 Z E D C B A gnd gnd vdd vdd
**PMOS current injection
Icharge 0 Z:F46 EXP (0 current_magnitude/3 rise_delay rise_time_constant fall_delay fall_time_constant)

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4_9

****** HS65_GS_AO212X4 : Glitched version 10 : glitch at Z:F56 ******

.SUBCKT HS65_GS_AO212X4_10 Z E D C B A gnd gnd vdd vdd
**PMOS current injection
Icharge 0 Z:F56 EXP (0 current_magnitude/3 rise_delay rise_time_constant fall_delay fall_time_constant)

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4_10

****** HS65_GS_AO212X4 : Glitched version 11 : glitch at net065:F38 ******

.SUBCKT HS65_GS_AO212X4_11 Z E D C B A gnd gnd vdd vdd
**NMOS current injection
Icharge net065:F38 0 EXP (0 current_magnitude rise_delay rise_time_constant fall_delay fall_time_constant)

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4_11

****** HS65_GS_AO212X4 : Glitched version 12 : glitch at net061:F26 ******

.SUBCKT HS65_GS_AO212X4_12 Z E D C B A gnd gnd vdd vdd
**NMOS current injection
Icharge net061:F26 0 EXP (0 current_magnitude rise_delay rise_time_constant fall_delay fall_time_constant)

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4_12

****** HS65_GS_AO212X4 : Glitched version 13 : glitch at net029:F30 ******

.SUBCKT HS65_GS_AO212X4_13 Z E D C B A gnd gnd vdd vdd
**NMOS current injection
Icharge net029:F30 0 EXP (0 current_magnitude rise_delay rise_time_constant fall_delay fall_time_constant)

*COMMENT Extracted with DK_cmos065lpgp_RF_7m4x0y2z_2V51V8@5.0.2@20070413.0 at 12:03 14 May 2007
Xld_D0 gnd vdd DNWPS AREA=3.504 PJ=7.72
MMM0 net044:F64 E:F63 net040:F62 vdd PSVTGP L=0.06u W=0.51u ad=0.051p as=0.109167p lpe=3 ngcon=1 nrd=0.215686 nrs=0.41971 pd=0.2u po2act=0.336651 ps=1.34u sca=9.53146 scb=0.0101069 scc=0.000839115
MMM1 net029:F50 C:F51 net044:F52 vdd PSVTGP AD=0.0765p AS=0.1071p L=0.06u NRD=0.313725 NRS=0.235294 PD=0.3u PS=0.93u W=0.51u lpe=3 ngcon=1 po2act=0.342878 sca=9.53197 scb=0.0101069 scc=0.000839115
MMM10 net029:F42 B:F43 net065:F44 gnd NSVTGP AD=0.05115p AS=0.02015p L=0.06u NRD=0.177419 NRS=0.209677 PD=0.64u PS=0.13u W=0.31u lpe=3 ngcon=1 po2act=0.267407 sca=2.56233 scb=0.000870205 scc=1.93523e-06
MMM11 net029:F36 E:F35 gnd gnd NSVTGP L=0.06u W=0.2u ad=0.0240784p as=0.0259804p lpe=3 ngcon=1 nrd=0.35 nrs=0.0826531 pd=0.223529u po2act=0.775155 ps=0.227451u sca=2.86219 scb=0.00118863 scc=2.93513e-06
MMM2 net029:F60 D:F59 net044:F58 vdd PSVTGP L=0.06u W=0.51u ad=0.0765p as=0.051p lpe=3 ngcon=1 nrd=0.509804 nrs=0.215686 pd=0.3u po2act=0.553309 ps=0.2u sca=9.53143 scb=0.0101069 scc=0.000839115
MMM3 Z:F24 net029:F23 gnd gnd NSVTGP L=0.06u W=0.39u ad=0.0663p as=0.0468557p lpe=3 ngcon=1 nrd=0.307692 nrs=0.358974 pd=0.73u po2act=0.251217 ps=0.300857u sca=2.92667 scb=0.00139386 scc=6.60165e-06
MMM4 net040:F70 B:F71 vdd vdd PSVTGP AD=0.109167p AS=0.051p L=0.06u NRD=0.41971 NRS=0.215686 PD=1.34u PS=0.2u W=0.51u lpe=3 ngcon=1 po2act=0.227263 sca=2.76163 scb=0.00145073 scc=9.47451e-06
MMM5 net040:F68 A:F67 vdd vdd PSVTGP L=0.06u W=0.51u ad=0.109167p as=0.051p lpe=3 ngcon=1 nrd=0.41971 nrs=0.215686 pd=1.34u po2act=0.300468 ps=0.2u sca=2.76088 scb=0.00145073 scc=9.47451e-06
MMM6 Z:F46 net029:F47 vdd vdd PSVTGP AD=0.0454545p AS=0.04125p L=0.06u NRD=1.37778 NRS=0.22 PD=0.381818u PS=0.58u W=0.25u lpe=3 ngcon=1 po2act=0.254897 sca=1.1443 scb=1.64443e-05 scc=3.54779e-10
MMM6@2 Z:F56 net029:F55 vdd vdd PSVTGP L=0.06u W=0.3u ad=0.0545455p as=0.0615p lpe=3 ngcon=1 nrd=0.0911157 nrs=0.216667 pd=0.458182u po2act=0.276956 ps=0.71u sca=1.1763 scb=2.24363e-05 scc=7.69694e-10
MMM7 net065:F38 A:F39 gnd gnd NSVTGP AD=0.02015p AS=0.0402696p L=0.06u NRD=0.209677 NRS=0.177419 PD=0.13u PS=0.352549u W=0.31u lpe=3 ngcon=1 po2act=0.37323 sca=2.56201 scb=0.000870205 scc=1.93523e-06
MMM8 net061:F26 C:F27 gnd gnd NSVTGP AD=0.02325p AS=0.0372443p L=0.06u NRD=0.241935 NRS=0.225806 PD=0.15u PS=0.239143u W=0.31u lpe=3 ngcon=1 po2act=0.533511 sca=2.56188 scb=0.000870205 scc=1.93523e-06
MMM9 net029:F30 D:F31 net061:F32 gnd NSVTGP AD=0.0373216p AS=0.02325p L=0.06u NRD=0.225806 NRS=0.241935 PD=0.346471u PS=0.15u W=0.31u lpe=3 ngcon=1 po2act=0.424318 sca=2.56172 scb=0.000870205 scc=1.93523e-06
R1 net065:F38 net065:F44 0.001
R10 D D:F6 0.001
R11 D:F59 D:F6 73.5984
R12 D:F59 D:F31 236.51
R13 D:F6 D:F31 331.193
R14 C C:F5 0.001
R15 C:F51 C:F27 225.329
R16 C:F51 C:F5 68.0437
R17 C:F5 C:F27 369.643
R18 E E:F7 0.001
R19 E:F63 E:F7 266.776
R2 net061:F26 net061:F32 0.001
R20 E:F63 E:F35 253.593
R21 E:F7 E:F35 85.3299
R22 B B:F4 0.001
R23 B:F71 B:F4 151.118
R24 B:F71 B:F43 500.572
R25 B:F4 B:F43 218.479
R26 A A:F3 0.001
R27 A:F67 A:F39 509.146
R28 A:F67 A:F3 150.639
R29 A:F3 A:F39 219.269
R3 gnd gnd 0.001
R30 Z Z:F8 0.001
R31 Z:F46 Z:F56 0.001
R32 Z:F46 Z:F8 37.7441
R33 Z:F8 Z:F24 39.4269
R34 net029:F55 net029:F47 143.75
R35 net029:F47 net029:F50 2320.39
R36 net029:F47 net029:F42 2464.11
R37 net029:F47 net029:F30 2394.27
R38 net029:F47 net029:F23 566.01
R39 net029:F50 net029:F60 0.001
R4 gnd gnd 0.001
R40 net029:F50 net029:F42 142.703
R41 net029:F50 net029:F30 138.659
R42 net029:F50 net029:F23 270.182
R43 net029:F23 net029:F42 286.916
R44 net029:F23 net029:F30 278.784
R45 net029:F30 net029:F42 131.338
R46 net029:F30 net029:F36 0.001
R47 net040:F68 net040:F70 0.001
R48 net040:F68 net040:F62 0.001
R49 vdd vdd 0.001
R5 gnd gnd 37.6143
R50 vdd vdd 0.001
R51 vdd vdd 0.001
R52 vdd vdd 0.001
R53 vdd vdd 0.001
R54 vdd vdd 0.001
R55 vdd vdd 0.001
R56 vdd vdd 0.001
R57 vdd vdd 37.6252
R58 vdd vdd 0.001
R59 vdd vdd 38.2613
R6 gnd gnd 37.721
R60 vdd vdd 37.8019
R61 vdd vdd 37.5
R62 vdd vdd 0.001
R63 gnd gnd 0.001
R64 gnd gnd 0.0256454
R65 gnd gnd 37.6257
R66 gnd gnd 0.001
R67 gnd gnd 0.001
R68 gnd gnd 0.001
R69 gnd gnd 0.001
R7 gnd gnd 0.001
R70 gnd gnd 0.001
R8 net044:F52 net044:F58 75.7472
R9 net044:F58 net044:F64 0.001
.ENDS HS65_GS_AO212X4_13

		**************************************** LIBRARAY INFORMATION ****************************************
 **** This Library contains 1 glitch free Subcircuits 
 **** This Library contains 13 glitch affected Subcircuits 
 **** Following are the details of these Subcircuits


**** SUBCIRCUIT		|VERSION COUNT
**-----------------------------------------
**** HS65_GS_AO212X4		|	13
************************************************************ END ************************************************************